magic
tech scmos
timestamp 1415052506
<< metal1 >>
rect 2342 3992 2354 4004
rect 1008 3980 1334 3992
rect 1346 3980 1805 3992
rect 1817 3980 2276 3992
rect 2288 3980 2746 3992
rect 2758 3980 3218 3992
rect 3230 3980 3992 3992
rect 1008 1020 1020 3980
rect 1028 3960 3972 3972
rect 1028 1040 1040 3960
rect 1342 3753 1350 3759
rect 1813 3757 1820 3763
rect 1334 3661 1342 3662
rect 1342 3653 1351 3659
rect 1813 3657 1819 3663
rect 1742 3493 1816 3497
rect 1763 3102 1821 3106
rect 1366 3081 1738 3085
rect 1836 3081 2209 3085
rect 1275 3074 1738 3078
rect 1838 3074 2680 3078
rect 1382 3067 1518 3071
rect 1889 3067 1977 3071
rect 2680 2603 2684 2607
rect 3960 1040 3972 3960
rect 1028 1028 1766 1040
rect 1778 1028 2237 1040
rect 2249 1028 2642 1040
rect 2654 1028 2708 1040
rect 2720 1028 3179 1040
rect 3191 1028 3650 1040
rect 3662 1028 3972 1040
rect 3980 1020 3992 3980
rect 1008 1008 3992 1020
<< m2contact >>
rect 1334 3980 1346 3992
rect 1805 3980 1817 3992
rect 2276 3980 2288 3992
rect 2746 3980 2758 3992
rect 3218 3980 3230 3992
rect 1334 3753 1342 3761
rect 1805 3757 1813 3765
rect 1334 3653 1342 3661
rect 1805 3657 1813 3665
rect 1777 3631 1781 3635
rect 2248 3631 2252 3635
rect 2719 3631 2723 3635
rect 3190 3631 3194 3635
rect 3661 3631 3665 3635
rect 1784 3501 1788 3505
rect 2255 3501 2259 3505
rect 2726 3501 2730 3505
rect 3197 3501 3201 3505
rect 3668 3501 3672 3505
rect 1738 3493 1742 3497
rect 1738 3181 1742 3185
rect 1738 3151 1742 3155
rect 1327 3116 1331 3120
rect 1798 3116 1802 3120
rect 2269 3116 2273 3120
rect 2740 3116 2744 3120
rect 3211 3116 3215 3120
rect 1759 3102 1763 3106
rect 1320 3095 1324 3099
rect 1791 3095 1795 3099
rect 2262 3095 2266 3099
rect 2733 3095 2737 3099
rect 3204 3095 3208 3099
rect 1758 3088 1762 3092
rect 1362 3081 1366 3085
rect 1738 3081 1742 3085
rect 1832 3081 1836 3085
rect 2209 3081 2213 3085
rect 1738 3074 1742 3078
rect 1834 3074 1838 3078
rect 2680 3074 2684 3078
rect 1378 3067 1382 3071
rect 1518 3067 1522 3071
rect 1885 3067 1889 3071
rect 1977 3067 1981 3071
rect 1777 3053 1781 3057
rect 2248 3053 2252 3057
rect 2719 3053 2723 3057
rect 3190 3053 3194 3057
rect 3661 3053 3665 3057
rect 1784 2923 1788 2927
rect 2255 2923 2259 2927
rect 2726 2923 2730 2927
rect 3197 2923 3201 2927
rect 3668 2923 3672 2927
rect 1362 2915 1366 2919
rect 1834 2915 1838 2919
rect 1738 2603 1742 2607
rect 2209 2603 2213 2607
rect 1327 2538 1331 2542
rect 1798 2538 1802 2542
rect 2269 2538 2273 2542
rect 2740 2538 2744 2542
rect 3211 2538 3215 2542
rect 1320 2517 1324 2521
rect 1791 2517 1795 2521
rect 2262 2517 2266 2521
rect 2733 2517 2737 2521
rect 3204 2517 3208 2521
rect 1777 2475 1781 2479
rect 2248 2475 2252 2479
rect 2719 2475 2723 2479
rect 3190 2475 3194 2479
rect 3661 2475 3665 2479
rect 1784 2345 1788 2349
rect 2255 2345 2259 2349
rect 2726 2345 2730 2349
rect 3197 2345 3201 2349
rect 3668 2345 3672 2349
rect 1327 1960 1331 1964
rect 1798 1960 1802 1964
rect 2269 1960 2273 1964
rect 2740 1960 2744 1964
rect 3211 1960 3215 1964
rect 1320 1939 1324 1943
rect 1791 1939 1795 1943
rect 2262 1939 2266 1943
rect 2733 1939 2737 1943
rect 3204 1939 3208 1943
rect 1777 1897 1781 1901
rect 2248 1897 2252 1901
rect 2719 1897 2723 1901
rect 3190 1897 3194 1901
rect 3661 1897 3665 1901
rect 1784 1767 1788 1771
rect 2255 1767 2259 1771
rect 2726 1767 2730 1771
rect 3197 1767 3201 1771
rect 3668 1767 3672 1771
rect 1327 1382 1331 1386
rect 1798 1382 1802 1386
rect 2269 1382 2273 1386
rect 2740 1382 2744 1386
rect 3211 1382 3215 1386
rect 1320 1361 1324 1365
rect 1791 1361 1795 1365
rect 2262 1361 2266 1365
rect 2733 1361 2737 1365
rect 3204 1361 3208 1365
rect 1766 1028 1778 1040
rect 2237 1028 2249 1040
rect 2642 1028 2654 1040
rect 2708 1028 2720 1040
rect 3179 1028 3191 1040
rect 3650 1028 3662 1040
<< metal2 >>
rect 1334 3761 1342 3980
rect 1334 3661 1342 3753
rect 1320 2521 1324 3095
rect 1320 1943 1324 2517
rect 1320 1365 1324 1939
rect 1327 2542 1331 3116
rect 1327 1964 1331 2538
rect 1327 1386 1331 1960
rect 1334 1496 1342 3653
rect 1805 3765 1813 3980
rect 1805 3665 1813 3757
rect 1738 3185 1742 3493
rect 1738 3085 1742 3151
rect 1759 3092 1763 3102
rect 1762 3088 1763 3092
rect 1362 2919 1366 3081
rect 1738 2607 1742 3074
rect 1766 1040 1774 3508
rect 1777 3057 1781 3631
rect 1777 2479 1781 3053
rect 1777 1901 1781 2475
rect 1784 2927 1788 3501
rect 1784 2349 1788 2923
rect 1784 1771 1788 2345
rect 1791 2521 1795 3095
rect 1791 1943 1795 2517
rect 1791 1365 1795 1939
rect 1798 2542 1802 3116
rect 1798 1964 1802 2538
rect 1798 1386 1802 1960
rect 1805 1496 1813 3657
rect 1832 3085 1836 3366
rect 1834 2919 1838 3074
rect 1885 3062 1889 3067
rect 2209 2607 2213 3081
rect 1977 2486 1981 2493
rect 2237 1040 2245 3508
rect 2248 3057 2252 3631
rect 2248 2479 2252 3053
rect 2248 1901 2252 2475
rect 2255 2927 2259 3501
rect 2255 2349 2259 2923
rect 2255 1771 2259 2345
rect 2262 2521 2266 3095
rect 2262 1943 2266 2517
rect 2262 1365 2266 1939
rect 2269 2542 2273 3116
rect 2269 1964 2273 2538
rect 2269 1386 2273 1960
rect 2276 1495 2284 3980
rect 2680 2603 2684 3074
rect 2708 1040 2716 3508
rect 2719 3057 2723 3631
rect 2719 2479 2723 3053
rect 2719 1901 2723 2475
rect 2726 2927 2730 3501
rect 2726 2349 2730 2923
rect 2726 1771 2730 2345
rect 2733 2521 2737 3095
rect 2733 1943 2737 2517
rect 2733 1365 2737 1939
rect 2740 2542 2744 3116
rect 2740 1964 2744 2538
rect 2740 1386 2744 1960
rect 2747 1495 2755 3980
rect 3179 1040 3187 3273
rect 3190 3057 3194 3631
rect 3190 2479 3194 3053
rect 3190 1901 3194 2475
rect 3197 2927 3201 3501
rect 3197 2349 3201 2923
rect 3197 1771 3201 2345
rect 3204 2521 3208 3095
rect 3204 1943 3208 2517
rect 3204 1365 3208 1939
rect 3211 2542 3215 3116
rect 3211 1964 3215 2538
rect 3211 1386 3215 1960
rect 3218 1495 3226 3980
rect 3650 1405 3658 3508
rect 3661 3057 3665 3631
rect 3661 2479 3665 3053
rect 3661 1901 3665 2475
rect 3668 2927 3672 3501
rect 3668 2349 3672 2923
rect 3668 1771 3672 2345
rect 3650 1040 3658 1398
rect 2642 1000 2654 1028
rect 2708 1027 2716 1028
rect 3179 1027 3187 1028
rect 2602 996 2698 1000
rect 2620 994 2634 996
use DMUX  DMUX_0
timestamp 1414996929
transform 1 0 1358 0 1 3650
box -19 3 78 111
use MUX2X1  MUX2X1_0
timestamp 1414990262
transform 1 0 1815 0 1 3660
box -5 -3 53 105
use PLU  PLU_0
array 0 4 471 0 3 578
timestamp 1414992301
transform 1 0 1326 0 1 1377
box -9 -40 462 538
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1415033039
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
