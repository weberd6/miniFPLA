magic
tech scmos
timestamp 1416164212
<< metal1 >>
rect 2342 3992 2354 4004
rect 1008 3980 1309 3992
rect 1321 3980 1805 3992
rect 1817 3980 1910 3992
rect 1922 3980 2276 3992
rect 2288 3980 2743 3992
rect 2755 3980 2809 3992
rect 2821 3980 3218 3992
rect 3230 3989 3992 3992
rect 3230 3980 3980 3989
rect 1008 3421 1020 3980
rect 1008 3121 1020 3409
rect 1008 2822 1020 3109
rect 1008 2521 1020 2810
rect 1008 1921 1020 2509
rect 1008 1622 1020 1909
rect 1008 1322 1020 1610
rect 1008 1020 1020 1310
rect 1028 3960 1043 3972
rect 1055 3960 1353 3972
rect 1365 3960 1556 3972
rect 1568 3960 1610 3972
rect 1622 3960 2156 3972
rect 2554 3960 3055 3972
rect 3067 3960 3143 3972
rect 3155 3960 3409 3972
rect 3421 3960 3710 3972
rect 3722 3960 3972 3972
rect 1028 3754 1040 3960
rect 1782 3952 1859 3957
rect 3127 3953 3359 3957
rect 3590 3952 3938 3957
rect 3556 3769 3659 3773
rect 1872 3761 1946 3765
rect 2656 3761 2761 3765
rect 2814 3761 2846 3765
rect 3134 3762 3771 3766
rect 1250 3754 1818 3758
rect 1822 3754 2269 3758
rect 2273 3754 2659 3758
rect 2663 3754 2760 3758
rect 2764 3754 3130 3758
rect 1326 3745 1334 3751
rect 1813 3745 1820 3751
rect 2739 3745 2747 3751
rect 2755 3745 2766 3751
rect 3208 3745 3218 3751
rect 3226 3745 3554 3751
rect 3960 3744 3972 3960
rect 1028 3667 1040 3742
rect 1318 3714 1363 3718
rect 3202 3714 3248 3718
rect 3729 3686 3952 3690
rect 1851 3681 1864 3685
rect 2793 3681 2806 3685
rect 1239 3671 1250 3675
rect 1331 3669 1378 3673
rect 1860 3671 1864 3681
rect 2802 3671 2806 3681
rect 3215 3669 3262 3673
rect 2735 3666 2740 3667
rect 2324 3661 2652 3665
rect 2735 3664 2736 3666
rect 1354 3656 1438 3660
rect 1028 3368 1040 3655
rect 1882 3654 2209 3658
rect 2309 3654 2652 3658
rect 2824 3654 3097 3658
rect 1326 3645 1766 3651
rect 1774 3645 1814 3651
rect 1876 3645 2661 3651
rect 2739 3645 2770 3651
rect 2818 3645 3551 3651
rect 1330 3638 1356 3642
rect 1759 3638 1821 3642
rect 2230 3638 2300 3642
rect 2701 3638 2764 3642
rect 3172 3638 3234 3642
rect 1758 3631 1777 3635
rect 1781 3631 2248 3635
rect 2252 3631 2719 3635
rect 2723 3631 3190 3635
rect 3194 3631 3595 3635
rect 3599 3631 3661 3635
rect 1048 3627 1350 3631
rect 3101 3624 3151 3628
rect 1326 3608 1350 3614
rect 3673 3606 3952 3611
rect 1750 3548 1754 3552
rect 1224 3541 1235 3545
rect 1239 3541 1250 3545
rect 1327 3508 1346 3514
rect 1232 3501 1242 3505
rect 1742 3493 1838 3497
rect 2684 3493 2758 3497
rect 3960 3445 3972 3732
rect 1584 3369 1592 3373
rect 2057 3369 2063 3373
rect 2513 3369 2534 3373
rect 2984 3369 3005 3373
rect 3455 3369 3475 3373
rect 1324 3362 1354 3366
rect 1836 3362 1852 3366
rect 2213 3362 2287 3366
rect 3155 3362 3229 3366
rect 1028 3068 1040 3356
rect 3768 3349 3951 3354
rect 3626 3239 3683 3243
rect 3643 3223 3680 3229
rect 3705 3159 3721 3163
rect 3717 3150 3721 3159
rect 3960 3144 3972 3433
rect 3648 3123 3684 3129
rect 3551 3116 3585 3120
rect 3679 3116 3771 3120
rect 3581 3113 3585 3116
rect 3581 3109 3764 3113
rect 1317 3102 1350 3106
rect 1763 3102 1821 3106
rect 2234 3102 2292 3106
rect 2705 3102 2763 3106
rect 3176 3102 3233 3106
rect 3644 3088 3707 3092
rect 1292 3081 1355 3085
rect 1366 3081 1738 3085
rect 1836 3081 2209 3085
rect 2310 3081 2680 3085
rect 2779 3081 3151 3085
rect 3252 3081 3622 3085
rect 1268 3074 1738 3078
rect 1838 3074 2680 3078
rect 2781 3074 3622 3078
rect 1048 3067 1362 3071
rect 1382 3067 1518 3071
rect 1614 3067 1875 3071
rect 1889 3067 1977 3071
rect 2085 3067 2299 3071
rect 2324 3067 2460 3071
rect 2556 3067 2819 3071
rect 2831 3067 2919 3071
rect 3027 3067 3239 3071
rect 3266 3067 3402 3071
rect 1621 3060 1764 3064
rect 2093 3060 2235 3064
rect 2564 3060 2706 3064
rect 3034 3060 3177 3064
rect 3494 3060 3597 3064
rect 1028 2768 1040 3056
rect 3566 3046 3643 3050
rect 3730 3049 3952 3054
rect 1312 3030 1336 3036
rect 1224 2976 1260 2980
rect 1288 2966 1302 2970
rect 1298 2959 1302 2966
rect 1314 2930 1352 2936
rect 1048 2846 1305 2851
rect 3960 2844 3972 3132
rect 1571 2791 1592 2795
rect 2042 2791 2063 2795
rect 2513 2791 2534 2795
rect 2984 2791 3005 2795
rect 3455 2791 3476 2795
rect 3960 2791 3972 2832
rect 1028 2255 1040 2756
rect 3684 2654 3771 2658
rect 3645 2645 3686 2651
rect 3756 2611 3764 2614
rect 3650 2545 3680 2551
rect 3680 2536 3952 2541
rect 1764 2517 1788 2521
rect 2235 2517 2259 2521
rect 2706 2517 2730 2521
rect 3177 2517 3201 2521
rect 3647 2517 3753 2521
rect 1784 2510 1788 2517
rect 2255 2510 2259 2517
rect 2726 2510 2730 2517
rect 3197 2510 3201 2517
rect 1048 2503 1362 2507
rect 1366 2503 2209 2507
rect 2308 2503 3151 2507
rect 3250 2503 3764 2507
rect 1366 2496 1738 2500
rect 1837 2496 2209 2500
rect 2310 2496 2680 2500
rect 2779 2496 3151 2500
rect 3252 2496 3622 2500
rect 1382 2489 1518 2493
rect 1889 2489 1977 2493
rect 2324 2489 2460 2493
rect 2831 2489 2919 2493
rect 3266 2489 3402 2493
rect 3420 2489 3952 2493
rect 1317 2482 1354 2486
rect 1763 2482 1821 2486
rect 2234 2482 2300 2486
rect 2705 2482 2774 2486
rect 3176 2482 3234 2486
rect 1313 2452 1349 2458
rect 1224 2383 1234 2387
rect 1306 2372 1311 2374
rect 1306 2371 1307 2372
rect 1313 2352 1351 2358
rect 1048 2345 1229 2349
rect 1742 2337 1816 2341
rect 2684 2337 2758 2341
rect 1028 2167 1040 2243
rect 3960 2245 3972 2779
rect 1571 2213 1592 2217
rect 2042 2213 2063 2217
rect 2513 2213 2534 2217
rect 2984 2213 3005 2217
rect 3455 2213 3476 2217
rect 1311 2206 1356 2210
rect 2213 2206 2287 2210
rect 3155 2206 3229 2210
rect 1028 1867 1040 2155
rect 3730 2149 3952 2154
rect 3626 2083 3683 2087
rect 3645 2067 3676 2073
rect 3707 2003 3721 2007
rect 3717 1993 3721 2003
rect 3650 1967 3676 1973
rect 3679 1960 3771 1964
rect 1317 1946 1350 1950
rect 1763 1946 1821 1950
rect 2234 1946 2291 1950
rect 2705 1946 2763 1950
rect 3176 1946 3234 1950
rect 3960 1944 3972 2233
rect 3643 1932 3707 1936
rect 1366 1925 1738 1929
rect 1837 1925 2209 1929
rect 2309 1925 2680 1929
rect 2779 1925 3151 1929
rect 3252 1925 3622 1929
rect 1267 1918 1738 1922
rect 1839 1918 2680 1922
rect 2781 1918 3622 1922
rect 1291 1911 1355 1915
rect 1382 1911 1518 1915
rect 1614 1911 1878 1915
rect 1889 1911 1977 1915
rect 2085 1911 2297 1915
rect 2324 1911 2460 1915
rect 2556 1911 2820 1915
rect 2831 1911 2919 1915
rect 3027 1911 3241 1915
rect 3266 1911 3402 1915
rect 1621 1904 1764 1908
rect 2093 1904 2235 1908
rect 2563 1904 2706 1908
rect 3035 1904 3177 1908
rect 3494 1904 3597 1908
rect 1048 1896 1362 1900
rect 2191 1890 2248 1894
rect 3565 1890 3643 1894
rect 1313 1874 1349 1880
rect 1028 1568 1040 1855
rect 1224 1820 1259 1824
rect 1287 1810 1301 1814
rect 1297 1802 1301 1810
rect 1311 1774 1352 1780
rect 1048 1646 1304 1651
rect 3960 1644 3972 1932
rect 1571 1635 1592 1639
rect 2042 1635 2063 1639
rect 2513 1635 2534 1639
rect 2984 1635 3004 1639
rect 3455 1635 3476 1639
rect 1028 1040 1040 1556
rect 3960 1591 3972 1632
rect 3684 1498 3771 1502
rect 3645 1489 3682 1495
rect 3756 1453 3764 1456
rect 3650 1389 3681 1395
rect 1781 1382 1798 1386
rect 1802 1382 1806 1386
rect 3680 1368 3951 1373
rect 1764 1361 1788 1365
rect 2235 1361 2259 1365
rect 2705 1361 2730 1365
rect 3177 1361 3201 1365
rect 3647 1361 3757 1365
rect 1317 1354 1319 1358
rect 1784 1354 1788 1361
rect 2255 1354 2259 1361
rect 2726 1354 2730 1361
rect 3197 1354 3201 1361
rect 1350 1347 1362 1351
rect 1366 1347 2209 1351
rect 2308 1347 3151 1351
rect 3250 1347 3764 1351
rect 1342 1338 1709 1344
rect 1760 1338 1796 1344
rect 1876 1338 2654 1344
rect 2705 1338 3098 1344
rect 3175 1338 3636 1344
rect 3649 1338 3714 1344
rect 1522 1331 1698 1335
rect 1882 1331 1977 1335
rect 1993 1330 2248 1334
rect 2464 1331 2639 1335
rect 2923 1330 3081 1334
rect 3406 1331 3584 1335
rect 1049 1323 1690 1327
rect 2779 1323 3088 1327
rect 1742 1274 1755 1278
rect 2680 1274 2697 1278
rect 3624 1274 3639 1278
rect 1751 1264 1755 1274
rect 2693 1265 2697 1274
rect 3635 1265 3639 1274
rect 3717 1268 3952 1272
rect 1761 1238 1766 1244
rect 1774 1238 1799 1244
rect 3173 1238 3179 1244
rect 3658 1238 3706 1244
rect 1702 1231 1741 1235
rect 1755 1231 1989 1235
rect 2643 1231 2682 1235
rect 3085 1231 3172 1235
rect 3588 1231 3625 1235
rect 1224 1224 1709 1228
rect 1713 1224 1798 1228
rect 2654 1224 3095 1228
rect 3099 1224 3593 1228
rect 3597 1224 3771 1228
rect 1210 1217 1320 1221
rect 1324 1217 1889 1221
rect 1893 1217 2262 1221
rect 2266 1217 2733 1221
rect 2737 1217 3204 1221
rect 1264 1210 1327 1214
rect 1331 1210 1777 1214
rect 1781 1210 2269 1214
rect 2273 1210 2740 1214
rect 2744 1210 3211 1214
rect 1694 1203 1751 1207
rect 1788 1202 2255 1206
rect 2259 1202 2459 1206
rect 2464 1202 2726 1206
rect 2730 1202 3197 1206
rect 3201 1202 3668 1206
rect 3960 1065 3972 1579
rect 1651 1043 1758 1048
rect 1796 1043 2159 1048
rect 2705 1043 2846 1048
rect 3093 1043 3359 1048
rect 3451 1043 3642 1048
rect 3960 1040 3972 1053
rect 1028 1028 1043 1040
rect 1055 1028 1555 1040
rect 1567 1028 1766 1040
rect 1778 1028 1856 1040
rect 1868 1028 1910 1040
rect 1922 1028 2210 1040
rect 2222 1028 2237 1040
rect 2249 1028 2708 1040
rect 2720 1028 3055 1040
rect 3067 1028 3110 1040
rect 3122 1028 3179 1040
rect 3191 1028 3648 1040
rect 3660 1028 3710 1040
rect 3722 1028 3972 1040
rect 3980 3690 3992 3977
rect 3980 3390 3992 3678
rect 3980 3089 3992 3378
rect 3980 2491 3992 3077
rect 3980 2191 3992 2479
rect 3980 1890 3992 2179
rect 3980 1858 3992 1878
rect 3980 1290 3992 1846
rect 1008 1008 1310 1020
rect 1322 1008 1610 1020
rect 2641 993 2653 1028
rect 3980 1020 3992 1278
rect 2821 1008 3409 1020
rect 3421 1008 3992 1020
<< m2contact >>
rect 1309 3980 1321 3992
rect 1805 3980 1817 3992
rect 1910 3980 1922 3992
rect 2276 3980 2288 3992
rect 2743 3980 2755 3992
rect 2809 3980 2821 3992
rect 3218 3980 3230 3992
rect 3980 3977 3992 3989
rect 1008 3409 1020 3421
rect 1008 3109 1020 3121
rect 1008 2810 1020 2822
rect 1008 2509 1020 2521
rect 1008 1909 1020 1921
rect 1008 1610 1020 1622
rect 1008 1310 1020 1322
rect 1043 3960 1055 3972
rect 1353 3960 1365 3972
rect 1556 3960 1568 3972
rect 1610 3960 1622 3972
rect 2156 3960 2168 3972
rect 2542 3960 2554 3972
rect 3055 3960 3067 3972
rect 3143 3960 3155 3972
rect 3409 3960 3421 3972
rect 3710 3960 3722 3972
rect 1777 3952 1782 3957
rect 1859 3952 1864 3957
rect 3123 3953 3127 3957
rect 3359 3952 3364 3957
rect 3585 3952 3590 3957
rect 3938 3952 3943 3957
rect 3552 3769 3556 3773
rect 3659 3769 3664 3774
rect 1868 3761 1872 3765
rect 1946 3761 1951 3766
rect 2652 3761 2656 3765
rect 2761 3761 2766 3766
rect 2810 3761 2814 3765
rect 2846 3761 2851 3766
rect 3130 3762 3134 3766
rect 3771 3762 3775 3766
rect 1246 3754 1250 3758
rect 1818 3754 1822 3758
rect 2269 3754 2273 3758
rect 2659 3754 2663 3758
rect 2760 3754 2764 3758
rect 3130 3754 3134 3758
rect 1028 3742 1040 3754
rect 1334 3743 1342 3751
rect 1805 3743 1813 3751
rect 2276 3743 2284 3751
rect 2747 3743 2755 3751
rect 3218 3743 3226 3751
rect 3960 3732 3972 3744
rect 1363 3714 1367 3718
rect 1868 3715 1872 3719
rect 2810 3713 2814 3717
rect 3248 3714 3252 3718
rect 1818 3691 1822 3695
rect 1826 3691 1830 3695
rect 1850 3691 1854 3695
rect 2269 3691 2273 3695
rect 2760 3691 2764 3695
rect 2768 3691 2772 3695
rect 2792 3691 2796 3695
rect 3552 3691 3556 3695
rect 3585 3691 3589 3695
rect 3595 3691 3599 3695
rect 3952 3686 3957 3691
rect 2253 3681 2257 3685
rect 3668 3681 3672 3685
rect 1235 3671 1239 3675
rect 1327 3669 1331 3673
rect 1378 3669 1382 3673
rect 2245 3671 2249 3675
rect 3211 3669 3215 3673
rect 3262 3669 3266 3673
rect 1028 3655 1040 3667
rect 2320 3661 2324 3665
rect 2652 3661 2656 3665
rect 2736 3662 2740 3666
rect 1350 3656 1354 3660
rect 1438 3656 1442 3660
rect 1878 3654 1882 3658
rect 2209 3654 2213 3658
rect 2305 3654 2309 3658
rect 2652 3654 2656 3658
rect 2820 3654 2824 3658
rect 3097 3654 3101 3658
rect 1766 3645 1774 3653
rect 1326 3638 1330 3642
rect 1777 3631 1781 3635
rect 2248 3631 2252 3635
rect 2719 3631 2723 3635
rect 3190 3631 3194 3635
rect 3595 3631 3599 3635
rect 3661 3631 3665 3635
rect 1043 3626 1048 3631
rect 1350 3627 1354 3631
rect 3097 3624 3101 3628
rect 3151 3624 3155 3628
rect 3668 3606 3673 3611
rect 3952 3606 3957 3611
rect 1220 3541 1224 3545
rect 1235 3541 1239 3545
rect 1320 3525 1324 3529
rect 1227 3501 1232 3506
rect 1242 3501 1246 3505
rect 1784 3501 1788 3505
rect 2255 3501 2259 3505
rect 2726 3501 2730 3505
rect 3197 3501 3201 3505
rect 3668 3501 3672 3505
rect 1363 3493 1367 3497
rect 1738 3493 1742 3497
rect 2305 3493 2309 3497
rect 2680 3493 2684 3497
rect 3248 3493 3252 3497
rect 3960 3433 3972 3445
rect 1028 3356 1040 3368
rect 1320 3362 1324 3366
rect 1832 3362 1836 3366
rect 2209 3362 2213 3366
rect 2775 3362 2779 3366
rect 3151 3362 3155 3366
rect 3763 3349 3768 3354
rect 3951 3349 3956 3354
rect 3622 3239 3626 3243
rect 3683 3239 3687 3243
rect 1738 3181 1742 3185
rect 2209 3181 2213 3185
rect 2680 3181 2684 3185
rect 3151 3181 3155 3185
rect 3622 3181 3626 3185
rect 3675 3169 3679 3173
rect 3683 3169 3687 3173
rect 3707 3169 3711 3173
rect 1738 3151 1742 3155
rect 2680 3151 2684 3155
rect 3622 3151 3626 3155
rect 3725 3154 3729 3158
rect 3960 3132 3972 3144
rect 1327 3116 1331 3120
rect 1798 3116 1802 3120
rect 2269 3116 2273 3120
rect 2740 3116 2744 3120
rect 3211 3116 3215 3120
rect 3675 3116 3679 3120
rect 3771 3116 3775 3120
rect 3764 3109 3768 3113
rect 1313 3102 1317 3106
rect 1759 3102 1763 3106
rect 2230 3102 2234 3106
rect 2701 3102 2705 3106
rect 3172 3102 3176 3106
rect 1320 3095 1324 3099
rect 1791 3095 1795 3099
rect 2262 3095 2266 3099
rect 2733 3095 2737 3099
rect 3204 3095 3208 3099
rect 1758 3088 1762 3092
rect 2230 3088 2234 3092
rect 2701 3088 2705 3092
rect 3172 3088 3176 3092
rect 3707 3088 3711 3092
rect 1288 3081 1292 3085
rect 1355 3081 1359 3085
rect 1362 3081 1366 3085
rect 1738 3081 1742 3085
rect 1832 3081 1836 3085
rect 2209 3081 2213 3085
rect 2306 3081 2310 3085
rect 2680 3081 2684 3085
rect 2775 3081 2779 3085
rect 3151 3081 3155 3085
rect 3248 3081 3252 3085
rect 3622 3081 3626 3085
rect 1264 3074 1268 3078
rect 1738 3074 1742 3078
rect 1834 3074 1838 3078
rect 2680 3074 2684 3078
rect 2777 3074 2781 3078
rect 3622 3074 3626 3078
rect 1028 3056 1040 3068
rect 1043 3067 1048 3072
rect 1362 3067 1366 3071
rect 1378 3067 1382 3071
rect 1518 3067 1522 3071
rect 1610 3067 1614 3071
rect 1875 3067 1879 3071
rect 1885 3067 1889 3071
rect 1977 3067 1981 3071
rect 2081 3067 2085 3071
rect 2299 3067 2303 3071
rect 2320 3067 2324 3071
rect 2460 3067 2464 3071
rect 2552 3067 2556 3071
rect 2819 3067 2823 3071
rect 2827 3067 2831 3071
rect 2919 3067 2923 3071
rect 3023 3067 3027 3071
rect 3239 3067 3243 3071
rect 3262 3067 3266 3071
rect 3402 3067 3406 3071
rect 1617 3060 1621 3064
rect 2089 3060 2093 3064
rect 2560 3060 2564 3064
rect 3030 3060 3034 3064
rect 3597 3060 3601 3064
rect 1777 3053 1781 3057
rect 2248 3053 2252 3057
rect 2719 3053 2723 3057
rect 3190 3053 3194 3057
rect 3661 3053 3665 3057
rect 3562 3046 3566 3050
rect 3643 3046 3647 3050
rect 3725 3049 3730 3054
rect 3952 3049 3957 3054
rect 1220 2976 1224 2980
rect 1264 2976 1268 2980
rect 1288 2976 1292 2980
rect 1306 2966 1310 2970
rect 1784 2923 1788 2927
rect 2255 2923 2259 2927
rect 2726 2923 2730 2927
rect 3197 2923 3201 2927
rect 3668 2923 3672 2927
rect 1362 2915 1366 2919
rect 1834 2915 1838 2919
rect 2306 2915 2310 2919
rect 2777 2915 2781 2919
rect 3248 2915 3252 2919
rect 1043 2846 1048 2851
rect 1305 2846 1310 2851
rect 3960 2832 3972 2844
rect 1362 2784 1366 2788
rect 1833 2784 1837 2788
rect 2304 2784 2308 2788
rect 2775 2784 2779 2788
rect 3246 2784 3250 2788
rect 1028 2756 1040 2768
rect 3960 2779 3972 2791
rect 3680 2654 3684 2658
rect 3771 2654 3775 2658
rect 3764 2610 3768 2614
rect 1738 2603 1742 2607
rect 2209 2603 2213 2607
rect 2680 2603 2684 2607
rect 3151 2603 3155 2607
rect 3622 2603 3626 2607
rect 1738 2573 1742 2577
rect 2209 2573 2213 2577
rect 2680 2573 2684 2577
rect 3151 2573 3155 2577
rect 3622 2573 3626 2577
rect 1327 2538 1331 2542
rect 1798 2538 1802 2542
rect 2269 2538 2273 2542
rect 2740 2538 2744 2542
rect 3211 2538 3215 2542
rect 3675 2536 3680 2541
rect 3952 2536 3957 2541
rect 1320 2517 1324 2521
rect 1791 2517 1795 2521
rect 2262 2517 2266 2521
rect 2733 2517 2737 2521
rect 3204 2517 3208 2521
rect 3753 2517 3757 2521
rect 1313 2510 1317 2514
rect 1043 2503 1048 2508
rect 1362 2503 1366 2507
rect 2209 2503 2213 2507
rect 2304 2503 2308 2507
rect 3151 2503 3155 2507
rect 3246 2503 3250 2507
rect 3764 2503 3768 2507
rect 1362 2496 1366 2500
rect 1738 2496 1742 2500
rect 1833 2496 1837 2500
rect 2209 2496 2213 2500
rect 2306 2496 2310 2500
rect 2680 2496 2684 2500
rect 2775 2496 2779 2500
rect 3151 2496 3155 2500
rect 3248 2496 3252 2500
rect 3622 2496 3626 2500
rect 1378 2489 1382 2493
rect 1518 2489 1522 2493
rect 1885 2489 1889 2493
rect 1977 2489 1981 2493
rect 2320 2489 2324 2493
rect 2460 2489 2464 2493
rect 2827 2489 2831 2493
rect 2919 2489 2923 2493
rect 3262 2489 3266 2493
rect 3402 2489 3406 2493
rect 3416 2489 3420 2493
rect 3952 2488 3957 2493
rect 1313 2482 1317 2486
rect 1777 2475 1781 2479
rect 2248 2475 2252 2479
rect 2719 2475 2723 2479
rect 3190 2475 3194 2479
rect 3661 2475 3665 2479
rect 1220 2383 1224 2387
rect 1307 2368 1311 2372
rect 1043 2345 1048 2350
rect 1229 2345 1233 2349
rect 1784 2345 1788 2349
rect 2255 2345 2259 2349
rect 2726 2345 2730 2349
rect 3197 2345 3201 2349
rect 3668 2345 3672 2349
rect 1362 2337 1366 2341
rect 1738 2337 1742 2341
rect 2306 2337 2310 2341
rect 2680 2337 2684 2341
rect 3248 2337 3252 2341
rect 1028 2243 1040 2255
rect 3960 2233 3972 2245
rect 1307 2206 1311 2210
rect 1833 2206 1837 2210
rect 2209 2206 2213 2210
rect 2775 2206 2779 2210
rect 3151 2206 3155 2210
rect 1028 2155 1040 2167
rect 3725 2149 3730 2154
rect 3952 2149 3957 2154
rect 3622 2083 3626 2087
rect 3683 2083 3687 2087
rect 1738 2025 1742 2029
rect 2209 2025 2213 2029
rect 2680 2025 2684 2029
rect 3151 2025 3155 2029
rect 3622 2025 3626 2029
rect 3675 2013 3679 2017
rect 3683 2013 3687 2017
rect 3707 2013 3711 2017
rect 3725 2007 3729 2011
rect 1738 1995 1742 1999
rect 2209 1995 2213 1999
rect 2680 1995 2684 1999
rect 3622 1995 3626 1999
rect 1327 1960 1331 1964
rect 1798 1960 1802 1964
rect 2269 1960 2273 1964
rect 2740 1960 2744 1964
rect 3211 1960 3215 1964
rect 3675 1960 3679 1964
rect 3771 1960 3775 1964
rect 1313 1946 1317 1950
rect 1759 1946 1763 1950
rect 2230 1946 2234 1950
rect 2701 1946 2705 1950
rect 3172 1946 3176 1950
rect 1320 1939 1324 1943
rect 1791 1939 1795 1943
rect 2262 1939 2266 1943
rect 2733 1939 2737 1943
rect 3204 1939 3208 1943
rect 1759 1932 1763 1936
rect 2230 1932 2234 1936
rect 2701 1932 2705 1936
rect 3172 1932 3176 1936
rect 3707 1932 3711 1936
rect 3960 1932 3972 1944
rect 1362 1925 1366 1929
rect 1738 1925 1742 1929
rect 1833 1925 1837 1929
rect 2209 1925 2213 1929
rect 2305 1925 2309 1929
rect 2680 1925 2684 1929
rect 2775 1925 2779 1929
rect 3151 1925 3155 1929
rect 3248 1925 3252 1929
rect 3622 1925 3626 1929
rect 1263 1918 1267 1922
rect 1738 1918 1742 1922
rect 1835 1918 1839 1922
rect 2680 1918 2684 1922
rect 2777 1918 2781 1922
rect 3622 1918 3626 1922
rect 1287 1911 1291 1915
rect 1355 1911 1359 1915
rect 1378 1911 1382 1915
rect 1518 1911 1522 1915
rect 1610 1911 1614 1915
rect 1878 1911 1882 1915
rect 1885 1911 1889 1915
rect 1977 1911 1981 1915
rect 2081 1911 2085 1915
rect 2297 1911 2301 1915
rect 2320 1911 2324 1915
rect 2460 1911 2464 1915
rect 2552 1911 2556 1915
rect 2820 1911 2824 1915
rect 2827 1911 2831 1915
rect 2919 1911 2923 1915
rect 3023 1911 3027 1915
rect 3241 1911 3245 1915
rect 3262 1911 3266 1915
rect 3402 1911 3406 1915
rect 1617 1904 1621 1908
rect 2089 1904 2093 1908
rect 2559 1904 2563 1908
rect 3031 1904 3035 1908
rect 3597 1904 3601 1908
rect 1043 1896 1048 1901
rect 1362 1896 1366 1900
rect 1777 1897 1781 1901
rect 2248 1897 2252 1901
rect 2719 1897 2723 1901
rect 3190 1897 3194 1901
rect 3661 1897 3665 1901
rect 2187 1890 2191 1894
rect 2248 1890 2252 1894
rect 3561 1890 3565 1894
rect 3643 1890 3647 1894
rect 1028 1855 1040 1867
rect 1220 1820 1224 1824
rect 1263 1820 1267 1824
rect 1287 1820 1291 1824
rect 1305 1810 1309 1814
rect 1784 1767 1788 1771
rect 2255 1767 2259 1771
rect 2726 1767 2730 1771
rect 3197 1767 3201 1771
rect 3668 1767 3672 1771
rect 1362 1759 1366 1763
rect 1835 1759 1839 1763
rect 2305 1759 2309 1763
rect 2777 1759 2781 1763
rect 3248 1759 3252 1763
rect 1043 1646 1048 1651
rect 1304 1646 1309 1651
rect 3960 1632 3972 1644
rect 1362 1628 1366 1632
rect 1833 1628 1837 1632
rect 2304 1628 2308 1632
rect 2775 1628 2779 1632
rect 3246 1628 3250 1632
rect 1028 1556 1040 1568
rect 3960 1579 3972 1591
rect 3680 1498 3684 1502
rect 3771 1498 3775 1502
rect 3764 1452 3768 1456
rect 1738 1447 1742 1451
rect 2209 1447 2213 1451
rect 2680 1447 2684 1451
rect 3151 1447 3155 1451
rect 3622 1447 3626 1451
rect 1738 1417 1742 1421
rect 2209 1417 2213 1421
rect 2680 1417 2684 1421
rect 3151 1417 3155 1421
rect 3622 1417 3626 1421
rect 1327 1382 1331 1386
rect 1777 1382 1781 1386
rect 1798 1382 1802 1386
rect 2269 1382 2273 1386
rect 2740 1382 2744 1386
rect 3211 1382 3215 1386
rect 3675 1368 3680 1373
rect 3951 1368 3956 1373
rect 1320 1361 1324 1365
rect 1791 1361 1795 1365
rect 1889 1361 1893 1365
rect 2262 1361 2266 1365
rect 2733 1361 2737 1365
rect 3204 1361 3208 1365
rect 3757 1361 3761 1365
rect 1313 1354 1317 1358
rect 1346 1347 1350 1351
rect 1362 1347 1366 1351
rect 2209 1347 2213 1351
rect 2304 1347 2308 1351
rect 3151 1347 3155 1351
rect 3246 1347 3250 1351
rect 3764 1347 3768 1351
rect 1334 1336 1342 1344
rect 1518 1331 1522 1335
rect 1698 1331 1702 1335
rect 1878 1331 1882 1335
rect 1977 1331 1981 1335
rect 1989 1330 1993 1334
rect 2248 1330 2252 1334
rect 2460 1331 2464 1335
rect 2639 1331 2643 1335
rect 2919 1330 2923 1334
rect 3081 1330 3085 1334
rect 3402 1331 3406 1335
rect 3584 1331 3588 1335
rect 1043 1323 1049 1329
rect 1690 1323 1694 1327
rect 2775 1323 2779 1327
rect 3088 1323 3092 1327
rect 3167 1307 3171 1311
rect 1870 1303 1874 1307
rect 1709 1284 1713 1288
rect 1717 1284 1721 1288
rect 1741 1284 1745 1288
rect 2650 1284 2654 1288
rect 2658 1284 2662 1288
rect 2682 1284 2686 1288
rect 3593 1284 3597 1288
rect 3601 1284 3605 1288
rect 3625 1284 3629 1288
rect 1759 1274 1763 1278
rect 2701 1275 2705 1279
rect 1798 1264 1802 1268
rect 3095 1268 3099 1272
rect 3643 1270 3647 1274
rect 3705 1264 3709 1268
rect 3952 1267 3957 1272
rect 1766 1238 1774 1246
rect 2708 1236 2716 1244
rect 3179 1238 3187 1246
rect 3650 1238 3658 1246
rect 1698 1231 1702 1235
rect 1741 1231 1745 1235
rect 1751 1231 1755 1235
rect 1989 1231 1993 1235
rect 2639 1231 2643 1235
rect 2682 1231 2686 1235
rect 3081 1231 3085 1235
rect 3172 1231 3176 1235
rect 3584 1231 3588 1235
rect 3625 1231 3629 1235
rect 1220 1224 1224 1228
rect 1709 1224 1713 1228
rect 1798 1224 1802 1228
rect 2650 1224 2654 1228
rect 3095 1224 3099 1228
rect 3593 1224 3597 1228
rect 3771 1224 3775 1228
rect 1205 1217 1210 1222
rect 1320 1217 1324 1221
rect 1889 1217 1893 1221
rect 2262 1217 2266 1221
rect 2733 1217 2737 1221
rect 3204 1217 3208 1221
rect 1259 1209 1264 1214
rect 1327 1210 1331 1214
rect 1777 1210 1781 1214
rect 2269 1210 2273 1214
rect 2740 1210 2744 1214
rect 3211 1210 3215 1214
rect 1690 1203 1694 1207
rect 1751 1203 1755 1207
rect 1784 1202 1788 1206
rect 2255 1202 2259 1206
rect 2459 1202 2464 1207
rect 2726 1202 2730 1206
rect 3197 1202 3201 1206
rect 3668 1202 3672 1206
rect 3960 1053 3972 1065
rect 1646 1043 1651 1048
rect 1758 1043 1763 1048
rect 1791 1043 1796 1048
rect 2159 1043 2164 1048
rect 2700 1043 2705 1048
rect 2846 1043 2851 1048
rect 3088 1043 3093 1048
rect 3359 1043 3364 1048
rect 3446 1043 3451 1048
rect 3642 1043 3647 1048
rect 1043 1028 1055 1040
rect 1555 1028 1567 1040
rect 1766 1028 1778 1040
rect 1856 1028 1868 1040
rect 1910 1028 1922 1040
rect 2210 1028 2222 1040
rect 2237 1028 2249 1040
rect 2708 1028 2720 1040
rect 3055 1028 3067 1040
rect 3110 1028 3122 1040
rect 3179 1028 3191 1040
rect 3648 1028 3660 1040
rect 3710 1028 3722 1040
rect 3980 3678 3992 3690
rect 3980 3378 3992 3390
rect 3980 3077 3992 3089
rect 3980 2479 3992 2491
rect 3980 2179 3992 2191
rect 3980 1878 3992 1890
rect 3980 1846 3992 1858
rect 3980 1278 3992 1290
rect 1310 1008 1322 1020
rect 1610 1008 1622 1020
rect 2809 1008 2821 1020
rect 3409 1008 3421 1020
<< metal2 >>
rect 1011 3995 1020 4000
rect 1044 3995 1053 4000
rect 1011 3986 1053 3995
rect 1044 3972 1053 3986
rect 997 3959 1013 3964
rect 1008 3955 1013 3959
rect 1008 3950 1232 3955
rect 1000 3744 1028 3753
rect 1004 3720 1013 3744
rect 1000 3711 1013 3720
rect 1000 3657 1028 3666
rect 1043 3451 1048 3626
rect 1000 3446 1048 3451
rect 1000 3411 1008 3420
rect 1000 3357 1028 3366
rect 1000 3146 1048 3151
rect 1000 3111 1008 3120
rect 1043 3072 1048 3146
rect 1000 3057 1028 3066
rect 1220 2980 1224 3541
rect 1227 3506 1232 3950
rect 1259 3770 1264 4000
rect 1311 3992 1320 4000
rect 1344 3996 1353 4000
rect 1344 3987 1364 3996
rect 1311 3972 1319 3980
rect 1355 3972 1364 3987
rect 1557 3972 1566 4000
rect 1611 3995 1620 4000
rect 1644 3995 1653 4000
rect 1611 3986 1653 3995
rect 1611 3972 1620 3986
rect 1311 3964 1342 3972
rect 1236 3765 1264 3770
rect 1236 3691 1241 3765
rect 1246 3706 1250 3754
rect 1334 3751 1342 3964
rect 1235 3545 1239 3671
rect 1322 3669 1327 3673
rect 1242 3505 1246 3554
rect 1326 3532 1330 3638
rect 1320 3366 1324 3525
rect 1264 2980 1268 3074
rect 1288 2980 1292 3081
rect 1000 2846 1043 2851
rect 1000 2811 1008 2820
rect 1000 2757 1028 2766
rect 1000 2546 1048 2551
rect 1000 2511 1008 2520
rect 1043 2508 1048 2546
rect 996 2459 1048 2464
rect 1043 2350 1048 2459
rect 1220 2387 1224 2976
rect 1306 2851 1310 2966
rect 1313 2514 1317 3102
rect 1320 2521 1324 3095
rect 1000 2244 1028 2253
rect 1005 2220 1014 2244
rect 1000 2211 1014 2220
rect 1000 2157 1028 2166
rect 1000 1946 1048 1951
rect 1000 1911 1008 1920
rect 1043 1901 1048 1946
rect 1000 1857 1028 1866
rect 1220 1824 1224 2383
rect 1229 2349 1233 2398
rect 1313 2380 1317 2482
rect 1311 2376 1317 2380
rect 1307 2210 1311 2368
rect 1263 1824 1267 1918
rect 1287 1824 1291 1911
rect 1000 1646 1043 1651
rect 1000 1611 1008 1620
rect 1000 1557 1028 1566
rect 995 1347 1049 1351
rect 998 1345 1049 1347
rect 1043 1329 1049 1345
rect 1000 1311 1008 1320
rect 1000 1259 1210 1264
rect 1205 1222 1210 1259
rect 1220 1228 1224 1820
rect 1305 1651 1309 1810
rect 1313 1358 1317 1946
rect 1320 1943 1324 2517
rect 1320 1365 1324 1939
rect 1320 1221 1324 1361
rect 1327 2542 1331 3116
rect 1327 1964 1331 2538
rect 1327 1386 1331 1960
rect 1327 1214 1331 1382
rect 1334 1344 1342 3743
rect 1350 3631 1354 3656
rect 1363 3497 1367 3714
rect 1378 3638 1382 3669
rect 1438 3624 1442 3656
rect 1738 3185 1742 3493
rect 1532 3103 1536 3122
rect 1355 3092 1425 3096
rect 1355 3085 1359 3092
rect 1362 3071 1366 3081
rect 1362 2919 1366 3067
rect 1421 3060 1425 3092
rect 1738 3085 1742 3151
rect 1759 3092 1763 3102
rect 1762 3088 1763 3092
rect 1525 3078 1621 3082
rect 1525 3060 1529 3078
rect 1610 3060 1614 3067
rect 1617 3064 1621 3078
rect 1421 3056 1529 3060
rect 1362 2507 1366 2784
rect 1738 2607 1742 3074
rect 1738 2500 1742 2573
rect 1362 2341 1366 2496
rect 1738 2029 1742 2337
rect 1355 1936 1425 1940
rect 1355 1915 1359 1936
rect 1362 1900 1366 1925
rect 1421 1904 1425 1936
rect 1738 1929 1742 1995
rect 1759 1936 1763 1946
rect 1525 1922 1621 1926
rect 1525 1904 1529 1922
rect 1610 1904 1614 1911
rect 1617 1908 1621 1922
rect 1421 1900 1529 1904
rect 1362 1763 1366 1896
rect 1362 1351 1366 1628
rect 1738 1451 1742 1918
rect 1738 1379 1742 1417
rect 1350 1347 1351 1351
rect 1717 1375 1742 1379
rect 998 1044 1020 1053
rect 1011 1020 1020 1044
rect 1044 1020 1053 1028
rect 1000 1011 1053 1020
rect 1011 1000 1020 1011
rect 1044 1000 1053 1011
rect 1259 1000 1264 1209
rect 1311 1000 1320 1008
rect 1346 1000 1351 1347
rect 1518 1335 1522 1337
rect 1690 1207 1694 1323
rect 1698 1235 1702 1331
rect 1717 1288 1721 1375
rect 1709 1228 1713 1284
rect 1741 1235 1745 1284
rect 1751 1207 1755 1231
rect 1759 1048 1763 1274
rect 1766 1246 1774 3645
rect 1777 3635 1781 3952
rect 1777 3057 1781 3631
rect 1805 3751 1813 3980
rect 1859 3957 1864 4000
rect 1911 3992 1920 4000
rect 1946 3766 1951 4009
rect 2157 3972 2166 4000
rect 2511 3995 2520 4000
rect 2544 3995 2553 4000
rect 2511 3986 2553 3995
rect 1777 2479 1781 3053
rect 1777 1901 1781 2475
rect 1784 2927 1788 3501
rect 1784 2349 1788 2923
rect 1784 1771 1788 2345
rect 1557 1000 1566 1028
rect 1611 1000 1620 1008
rect 1646 1000 1651 1043
rect 1766 1040 1774 1238
rect 1777 1214 1781 1382
rect 1784 1206 1788 1767
rect 1791 2521 1795 3095
rect 1791 1943 1795 2517
rect 1791 1365 1795 1939
rect 1798 2542 1802 3116
rect 1798 1964 1802 2538
rect 1798 1386 1802 1960
rect 1805 1496 1813 3743
rect 1818 3695 1822 3754
rect 1868 3719 1872 3761
rect 2269 3695 2273 3754
rect 1854 3691 1889 3695
rect 2276 3751 2284 3980
rect 2544 3972 2553 3986
rect 1826 3658 1830 3691
rect 1826 3654 1878 3658
rect 1885 3629 1889 3691
rect 2209 3366 2213 3654
rect 2245 3644 2249 3671
rect 2253 3653 2257 3681
rect 2253 3649 2273 3653
rect 2245 3640 2266 3644
rect 1832 3085 1836 3362
rect 2209 3185 2213 3362
rect 2230 3092 2234 3102
rect 1875 3078 1897 3082
rect 1834 2919 1838 3074
rect 1875 3071 1879 3078
rect 1885 3062 1889 3067
rect 1893 3060 1897 3078
rect 1998 3078 2093 3082
rect 1998 3060 2002 3078
rect 2081 3060 2085 3067
rect 2089 3064 2093 3078
rect 1893 3056 2002 3060
rect 1833 2500 1837 2784
rect 2209 2607 2213 3081
rect 2209 2507 2213 2573
rect 1885 2482 1889 2489
rect 2209 2210 2213 2496
rect 1833 1929 1837 2206
rect 2209 2029 2213 2206
rect 2209 1954 2213 1995
rect 2187 1950 2213 1954
rect 1878 1922 1896 1926
rect 1835 1763 1839 1918
rect 1878 1915 1882 1922
rect 1885 1905 1889 1911
rect 1892 1904 1896 1922
rect 1997 1922 2093 1926
rect 1997 1904 2001 1922
rect 2081 1904 2085 1911
rect 2089 1908 2093 1922
rect 1892 1900 2001 1904
rect 2187 1894 2191 1950
rect 2230 1936 2234 1946
rect 1833 1347 1837 1628
rect 2209 1451 2213 1925
rect 1833 1343 1874 1347
rect 1870 1307 1874 1343
rect 1791 1048 1795 1288
rect 1878 1266 1882 1331
rect 1798 1228 1802 1264
rect 1871 1262 1882 1266
rect 1889 1221 1893 1361
rect 2209 1351 2213 1417
rect 1977 1335 1981 1341
rect 1989 1235 1993 1330
rect 1857 1000 1866 1028
rect 1911 1014 1920 1028
rect 1911 1005 1953 1014
rect 1911 1000 1920 1005
rect 1944 1000 1953 1005
rect 2159 1000 2164 1043
rect 2237 1040 2245 3508
rect 2248 3057 2252 3631
rect 2248 2479 2252 3053
rect 2248 1901 2252 2475
rect 2255 2927 2259 3501
rect 2255 2349 2259 2923
rect 2248 1334 2252 1890
rect 2255 1771 2259 2345
rect 2255 1206 2259 1767
rect 2262 3099 2266 3640
rect 2262 2521 2266 3095
rect 2262 1943 2266 2517
rect 2262 1365 2266 1939
rect 2262 1221 2266 1361
rect 2269 3120 2273 3649
rect 2269 2542 2273 3116
rect 2269 1964 2273 2538
rect 2269 1386 2273 1960
rect 2276 1495 2284 3743
rect 2652 3691 2656 3761
rect 2659 3706 2663 3754
rect 2747 3751 2755 3980
rect 2761 3766 2766 4009
rect 2811 3992 2820 4000
rect 2846 3766 2851 4000
rect 3057 3972 3066 4000
rect 3111 3994 3120 4000
rect 3144 3994 3153 4000
rect 3111 3985 3153 3994
rect 3144 3972 3153 3985
rect 2652 3669 2704 3673
rect 2652 3665 2656 3669
rect 2305 3497 2309 3654
rect 2320 3636 2324 3661
rect 2736 3658 2740 3662
rect 2656 3654 2740 3658
rect 2680 3185 2684 3493
rect 2299 3092 2372 3096
rect 2299 3071 2303 3092
rect 2306 2919 2310 3081
rect 2368 3060 2372 3092
rect 2680 3085 2684 3151
rect 2701 3092 2705 3102
rect 2468 3078 2564 3082
rect 2468 3060 2472 3078
rect 2552 3060 2556 3067
rect 2560 3064 2564 3078
rect 2368 3056 2472 3060
rect 2304 2507 2308 2784
rect 2680 2607 2684 3074
rect 2680 2500 2684 2573
rect 2306 2341 2310 2496
rect 2680 2029 2684 2337
rect 2297 1936 2367 1940
rect 2297 1915 2301 1936
rect 2305 1763 2309 1925
rect 2363 1904 2367 1936
rect 2680 1929 2684 1995
rect 2701 1936 2705 1946
rect 2467 1922 2563 1926
rect 2467 1904 2471 1922
rect 2552 1904 2556 1911
rect 2559 1908 2563 1922
rect 2363 1900 2471 1904
rect 2269 1214 2273 1382
rect 2304 1351 2308 1628
rect 2680 1451 2684 1918
rect 2680 1379 2684 1417
rect 2658 1375 2684 1379
rect 2460 1335 2464 1337
rect 2639 1235 2643 1331
rect 2658 1288 2662 1375
rect 2650 1228 2654 1284
rect 2682 1235 2686 1284
rect 2249 1028 2253 1040
rect 2211 1000 2220 1028
rect 2244 1000 2253 1028
rect 2459 1000 2464 1202
rect 2701 1048 2705 1275
rect 2708 1244 2716 3508
rect 2719 3057 2723 3631
rect 2719 2479 2723 3053
rect 2719 1901 2723 2475
rect 2726 2927 2730 3501
rect 2726 2349 2730 2923
rect 2708 1040 2716 1236
rect 2726 1771 2730 2345
rect 2726 1206 2730 1767
rect 2733 2521 2737 3095
rect 2733 1943 2737 2517
rect 2733 1365 2737 1939
rect 2733 1221 2737 1361
rect 2740 2542 2744 3116
rect 2740 1964 2744 2538
rect 2740 1386 2744 1960
rect 2747 1495 2755 3743
rect 2760 3695 2764 3754
rect 2810 3717 2814 3761
rect 2796 3691 2831 3695
rect 3123 3691 3127 3953
rect 3130 3758 3134 3762
rect 3130 3706 3134 3754
rect 3218 3751 3226 3980
rect 3359 3957 3364 4000
rect 3411 3996 3420 4000
rect 3444 3996 3453 4000
rect 3411 3987 3453 3996
rect 3411 3972 3420 3987
rect 2768 3658 2772 3691
rect 2768 3654 2820 3658
rect 2827 3638 2831 3691
rect 3207 3669 3211 3673
rect 3097 3628 3101 3654
rect 3151 3366 3155 3624
rect 2775 3085 2779 3362
rect 3151 3185 3155 3362
rect 3172 3092 3176 3102
rect 2819 3078 2843 3082
rect 2777 2919 2781 3074
rect 2819 3071 2823 3078
rect 2827 3060 2831 3067
rect 2839 3061 2843 3078
rect 2942 3078 3034 3082
rect 2942 3061 2946 3078
rect 2839 3057 2946 3061
rect 3023 3060 3027 3067
rect 3030 3064 3034 3078
rect 2775 2500 2779 2784
rect 3151 2607 3155 3081
rect 3151 2507 3155 2573
rect 2827 2482 2831 2489
rect 3151 2210 3155 2496
rect 2775 1929 2779 2206
rect 3151 2029 3155 2206
rect 3172 1936 3176 1946
rect 2820 1922 2838 1926
rect 2777 1763 2781 1918
rect 2820 1915 2824 1922
rect 2827 1898 2831 1911
rect 2834 1904 2838 1922
rect 2938 1922 3035 1926
rect 2938 1904 2942 1922
rect 3023 1904 3027 1911
rect 3031 1908 3035 1922
rect 2834 1900 2942 1904
rect 2740 1214 2744 1382
rect 2775 1327 2779 1628
rect 3151 1451 3155 1925
rect 3151 1351 3155 1417
rect 2919 1334 2923 1338
rect 3081 1235 3085 1330
rect 3088 1311 3092 1323
rect 3088 1307 3167 1311
rect 3088 1284 3093 1288
rect 3088 1048 3092 1284
rect 3095 1228 3099 1268
rect 3173 1262 3176 1266
rect 3172 1235 3176 1262
rect 3179 1246 3187 3273
rect 3190 3057 3194 3631
rect 3190 2479 3194 3053
rect 3190 1901 3194 2475
rect 3197 2927 3201 3501
rect 3197 2349 3201 2923
rect 2811 1000 2820 1008
rect 2846 1000 2851 1043
rect 3179 1040 3187 1238
rect 3197 1771 3201 2345
rect 3197 1206 3201 1767
rect 3204 2521 3208 3095
rect 3204 1943 3208 2517
rect 3204 1365 3208 1939
rect 3204 1221 3208 1361
rect 3211 2542 3215 3116
rect 3211 1964 3215 2538
rect 3211 1386 3215 1960
rect 3218 1495 3226 3743
rect 3248 3497 3252 3714
rect 3552 3695 3556 3769
rect 3585 3695 3589 3952
rect 3659 3774 3664 4000
rect 3711 3993 3720 4000
rect 3744 3993 3753 4000
rect 3711 3984 3753 3993
rect 3711 3972 3720 3984
rect 3959 3979 3964 4000
rect 3938 3974 3964 3979
rect 3992 3980 4000 3989
rect 3938 3957 3943 3974
rect 3952 3951 4000 3956
rect 3262 3645 3266 3669
rect 3595 3635 3599 3691
rect 3622 3185 3626 3239
rect 3239 3091 3315 3095
rect 3239 3071 3243 3091
rect 3248 2919 3252 3081
rect 3311 3060 3315 3091
rect 3409 3067 3566 3071
rect 3409 3060 3413 3067
rect 3311 3056 3413 3060
rect 3562 3050 3566 3067
rect 3597 3064 3601 3173
rect 3622 3085 3626 3151
rect 3246 2507 3250 2784
rect 3622 2607 3626 3074
rect 3643 3050 3647 3051
rect 3248 2341 3252 2496
rect 3416 2493 3420 2521
rect 3622 2500 3626 2573
rect 3622 2029 3626 2083
rect 3241 1936 3309 1940
rect 3241 1915 3245 1936
rect 3248 1763 3252 1925
rect 3305 1904 3309 1936
rect 3409 1911 3565 1915
rect 3409 1904 3413 1911
rect 3305 1900 3413 1904
rect 3561 1894 3565 1911
rect 3597 1908 3601 2017
rect 3622 1929 3626 1995
rect 3211 1214 3215 1382
rect 3246 1351 3250 1628
rect 3622 1451 3626 1918
rect 3622 1379 3626 1417
rect 3650 1405 3658 3508
rect 3661 3057 3665 3631
rect 3661 2479 3665 3053
rect 3661 1901 3665 2475
rect 3668 3611 3672 3681
rect 3668 3505 3672 3606
rect 3668 2927 3672 3501
rect 3683 3173 3687 3239
rect 3675 3120 3679 3169
rect 3707 3092 3711 3169
rect 3725 3158 3729 3163
rect 3725 3054 3729 3154
rect 3764 3113 3768 3349
rect 3771 3120 3775 3762
rect 3952 3691 3957 3951
rect 3972 3734 4000 3743
rect 3992 3680 4000 3689
rect 3952 3649 4000 3654
rect 3952 3611 3957 3649
rect 3972 3434 4000 3443
rect 3992 3380 4000 3389
rect 3956 3349 4000 3354
rect 3972 3134 4000 3143
rect 3668 2349 3672 2923
rect 3771 2658 3775 3116
rect 3992 3080 4000 3089
rect 3957 3049 4000 3054
rect 3972 2834 4000 2843
rect 3972 2780 4000 2789
rect 3986 2756 3995 2780
rect 3986 2747 4004 2756
rect 3680 2602 3684 2654
rect 3675 2541 3679 2595
rect 3753 2521 3757 2569
rect 3764 2507 3768 2610
rect 3668 1771 3672 2345
rect 3683 2017 3687 2083
rect 3675 1964 3679 2013
rect 3707 1936 3711 2013
rect 3725 2011 3729 2149
rect 3725 2003 3729 2007
rect 3771 1964 3775 2654
rect 3957 2536 4000 2541
rect 3952 2454 3957 2488
rect 3992 2480 4000 2489
rect 3952 2449 4000 2454
rect 3972 2234 4000 2243
rect 3992 2180 4000 2189
rect 3957 2149 4000 2154
rect 3601 1375 3626 1379
rect 3402 1335 3406 1340
rect 3584 1235 3588 1331
rect 3601 1288 3605 1375
rect 3593 1228 3597 1284
rect 3625 1235 3629 1284
rect 3643 1274 3647 1278
rect 3643 1048 3647 1270
rect 3057 1000 3066 1028
rect 3111 1014 3120 1028
rect 3111 1005 3153 1014
rect 3111 1000 3120 1005
rect 3144 1000 3153 1005
rect 3359 1000 3364 1043
rect 3650 1246 3658 1398
rect 3411 1000 3420 1008
rect 3446 1000 3451 1043
rect 3650 1040 3658 1238
rect 3668 1206 3672 1767
rect 3771 1502 3775 1960
rect 3972 1934 4000 1943
rect 3992 1880 4000 1889
rect 3992 1847 4000 1856
rect 3972 1634 4000 1643
rect 3972 1580 4000 1589
rect 3986 1556 3995 1580
rect 3986 1547 4000 1556
rect 3680 1450 3684 1498
rect 3675 1373 3679 1435
rect 3757 1365 3761 1417
rect 3764 1351 3768 1452
rect 3705 1049 3709 1264
rect 3771 1228 3775 1498
rect 3952 1341 3956 1368
rect 3952 1336 4000 1341
rect 3992 1280 4000 1289
rect 3952 1254 3957 1267
rect 3952 1249 4000 1254
rect 3972 1055 3984 1064
rect 3705 1043 3964 1049
rect 3650 1014 3659 1028
rect 3711 1014 3720 1028
rect 3650 1005 3666 1014
rect 3657 1000 3666 1005
rect 3711 1005 3753 1014
rect 3711 1000 3720 1005
rect 3744 1000 3753 1005
rect 3958 1000 3964 1043
rect 3975 1043 3984 1055
rect 3975 1034 4000 1043
rect 2602 996 2642 1000
rect 2654 996 2698 1000
rect 2620 994 2634 996
use DMUX  DMUX_0
timestamp 1416012586
transform 1 0 1254 0 1 3642
box -19 3 78 111
use MUX2X1  MUX2X1_5
timestamp 1414990262
transform 1 0 1816 0 1 3648
box -5 -3 53 105
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 1858 0 1 3648
box -9 -3 26 105
use OR2X1  OR2X1_0
timestamp 1053022145
transform 1 0 2243 0 1 3648
box -8 -3 40 105
use DMUX  DMUX_2
timestamp 1416012586
transform 1 0 2667 0 1 3642
box -19 3 78 111
use MUX2X1  MUX2X1_6
timestamp 1414990262
transform 1 0 2758 0 1 3648
box -5 -3 53 105
use INVX1  INVX1_1
timestamp 1053022145
transform 1 0 2800 0 1 3648
box -9 -3 26 105
use DMUX  DMUX_4
timestamp 1416012586
transform 1 0 3138 0 1 3642
box -19 3 78 111
use DFFPOSRL  DFFPOSRL_0
timestamp 1414990262
transform 1 0 3530 0 1 3382
box 16 256 205 376
use DMUX  DMUX_1
timestamp 1416012586
transform 1 0 1255 0 1 3505
box -19 3 78 111
use MUX2X1  MUX2X1_7
timestamp 1414990262
transform 1 0 3673 0 1 3126
box -5 -3 53 105
use INVX1  INVX1_7
timestamp 1053022145
transform 1 0 3715 0 1 3126
box -9 -3 26 105
use MUX2X1  MUX2X1_4
timestamp 1414990262
transform 1 0 1254 0 1 2933
box -5 -3 53 105
use INVX1  INVX1_2
timestamp 1053022145
transform 1 0 1296 0 1 2933
box -9 -3 26 105
use DMUX  DMUX_5
timestamp 1416012586
transform 1 0 3688 0 1 2542
box -19 3 78 111
use DMUX  DMUX_3
timestamp 1416012586
transform 1 0 1242 0 1 2349
box -19 3 78 111
use MUX2X1  MUX2X1_8
timestamp 1414990262
transform 1 0 3673 0 1 1970
box -5 -3 53 105
use INVX1  INVX1_8
timestamp 1053022145
transform 1 0 3715 0 1 1970
box -9 -3 26 105
use MUX2X1  MUX2X1_0
timestamp 1414990262
transform 1 0 1253 0 1 1777
box -5 -3 53 105
use INVX1  INVX1_3
timestamp 1053022145
transform 1 0 1295 0 1 1777
box -9 -3 26 105
use DMUX  DMUX_6
timestamp 1416012586
transform 1 0 3688 0 1 1386
box -19 3 78 111
use PLU  PLU_0
array 0 4 471 0 3 578
timestamp 1416027737
transform 1 0 1326 0 1 1377
box -9 -40 462 538
use MUX2X1  MUX2X1_1
timestamp 1414990262
transform 1 0 1707 0 1 1241
box -5 -3 53 105
use INVX1  INVX1_4
timestamp 1053022145
transform 1 0 1749 0 1 1241
box -9 -3 26 105
use DMUX  DMUX_7
timestamp 1416012586
transform 1 0 1806 0 1 1235
box -19 3 78 111
use MUX2X1  MUX2X1_2
timestamp 1414990262
transform 1 0 2648 0 1 1241
box -5 -3 53 105
use INVX1  INVX1_5
timestamp 1053022145
transform 1 0 2691 0 1 1241
box -9 -3 26 105
use DMUX  DMUX_8
timestamp 1416012586
transform 1 0 3103 0 1 1235
box -19 3 78 111
use MUX2X1  MUX2X1_3
timestamp 1414990262
transform 1 0 3591 0 1 1241
box -5 -3 53 105
use INVX1  INVX1_6
timestamp 1053022145
transform 1 0 3633 0 1 1241
box -9 -3 26 105
use INVX1  INVX1_9
timestamp 1053022145
transform 1 0 3703 0 1 1241
box -9 -3 26 105
<< labels >>
rlabel metal2 1261 3993 1261 3993 1 In0
rlabel metal2 1352 3993 1352 3993 1 Gnd_out
rlabel metal2 1861 3993 1861 3993 1 Reset
rlabel metal2 1948 3994 1948 3994 1 Out0
rlabel metal2 2763 3994 2763 3994 1 In1
rlabel metal2 2848 3994 2848 3994 1 Out1
rlabel metal2 3361 3994 3361 3994 1 In2
rlabel metal2 3661 3994 3661 3994 1 Load
rlabel metal2 3961 3994 3961 3994 1 D
rlabel metal2 3993 3952 3993 3952 1 Q
rlabel metal2 3994 3650 3994 3650 1 clk_out1
rlabel metal2 3994 3350 3994 3350 1 test_out
rlabel metal2 3994 3051 3994 3051 1 Out2
rlabel metal2 3994 2538 3994 2538 1 In3
rlabel metal2 3994 2450 3994 2450 1 Cfg_out
rlabel metal2 3994 2151 3994 2151 1 Out3
rlabel metal2 3994 1849 3994 1849 1 Vdd_out
rlabel metal2 3994 1337 3994 1337 1 In4
rlabel metal2 3994 1250 3994 1250 1 Inv_out
rlabel metal2 3960 1004 3960 1004 1 Inv_in
rlabel metal2 3448 1005 3448 1005 1 Out4
rlabel metal2 3360 1004 3360 1004 1 In5
rlabel metal2 2848 1005 2848 1005 1 Out5
rlabel metal2 2461 1007 2461 1007 1 Clk
rlabel metal2 2161 1004 2161 1004 1 In6
rlabel metal2 1648 1005 1648 1005 1 Out6
rlabel metal2 1261 1004 1261 1004 1 Test
rlabel metal2 1004 1260 1004 1260 1 Cfg
rlabel metal2 1005 1347 1005 1347 1 t11
rlabel metal2 1004 1647 1004 1647 1 Out7
rlabel metal2 1005 1947 1005 1947 1 t10
rlabel metal2 1005 2460 1005 2460 1 In7
rlabel metal2 1005 2547 1005 2547 1 t6
rlabel metal2 1005 3147 1005 3147 1 t0
rlabel metal2 1005 3447 1005 3447 1 Clk_out
rlabel metal2 1005 3960 1005 3960 1 In8
rlabel metal2 1005 2847 1005 2847 1 Out8
rlabel metal1 1351 3715 1351 3715 1 in0_D0
rlabel metal1 1353 3670 1353 3670 1 in0_D1
rlabel metal2 1328 3539 1328 3539 1 in8_D1
rlabel metal2 1322 3518 1322 3518 1 in8_D0
rlabel metal1 2346 3985 2346 3985 1 Vdd
rlabel metal1 2645 1033 2645 1033 1 Gnd
rlabel metal1 1788 3639 1788 3639 1 first_mux_shift
rlabel metal1 1783 2483 1783 2483 1 second_mux_shift
rlabel metal1 1751 3550 1751 3550 1 first_muxff_out
rlabel metal2 3685 3234 3685 3234 1 output4
rlabel metal2 2210 3237 2210 3237 1 output1
rlabel metal2 2682 3116 2682 3116 1 output2
rlabel metal2 3152 3238 3152 3238 1 output3
rlabel metal2 1739 2536 1739 2536 1 output5
rlabel metal2 2210 2540 2210 2540 1 output6
rlabel metal2 2681 2535 2681 2535 1 output7
rlabel metal2 3152 2538 3152 2538 1 output8
rlabel metal2 3623 2539 3623 2539 1 output9
rlabel metal2 1739 1959 1739 1959 1 output10
rlabel metal2 2210 1956 2210 1956 1 output11
rlabel metal2 2681 1953 2681 1953 1 output12
rlabel metal2 3153 2082 3153 2082 1 output13
rlabel metal2 3624 1961 3624 1961 1 output14
rlabel metal2 1738 1380 1738 1380 1 output15
rlabel metal2 2681 1381 2681 1381 1 output17
rlabel metal2 3152 1373 3152 1373 1 output18
rlabel metal2 3622 1377 3622 1377 1 output19
rlabel metal2 1740 3239 1740 3239 1 output0
rlabel metal2 1348 1004 1348 1004 1 t16
rlabel metal2 2210 1381 2210 1381 1 output16
rlabel metal2 2737 3656 2737 3656 1 in1_D0
rlabel metal1 2646 3663 2646 3663 1 in1_D1
rlabel metal1 3238 3715 3238 3715 1 in2_D0
rlabel metal1 3240 3670 3240 3670 1 in2_D1
rlabel metal2 3765 2590 3765 2590 1 in3_D0
rlabel metal2 3754 2526 3754 2526 1 in3_D1
rlabel metal2 3765 1423 3765 1423 1 in4_D0
rlabel metal1 3742 1362 3742 1362 1 in4_D1
rlabel metal1 3163 1233 3163 1233 1 in5_D1
rlabel metal1 3068 1325 3068 1325 1 in5_D0
rlabel metal2 1880 1269 1880 1269 1 in6_D1
rlabel metal2 1835 1353 1835 1353 1 in6_D0
rlabel metal2 1314 2382 1314 2382 1 in7_D1
rlabel metal2 1308 2347 1308 2347 1 in7_D0
rlabel metal1 1850 3363 1850 3363 1 inp1_1
rlabel metal1 2288 3756 2288 3756 1 Test_or_config
rlabel metal1 2059 3371 2059 3371 1 lut_out1
rlabel metal1 1586 3370 1586 3370 1 lut_out0
rlabel metal1 2528 3370 2528 3370 1 lut_out2
rlabel metal1 2998 3370 2998 3370 1 lut_out3
rlabel metal1 3470 3370 3470 3370 1 lut_out4
rlabel metal1 1585 2792 1585 2792 1 lut_out5
rlabel metal1 2056 2792 2056 2792 1 lut_out6
rlabel metal1 2528 2793 2528 2793 1 lut_out7
rlabel metal1 2998 2792 2998 2792 1 lut_out8
rlabel metal1 3469 2792 3469 2792 1 lut_out9
rlabel metal1 1585 2214 1585 2214 1 lut_out10
rlabel metal1 2057 2214 2057 2214 1 lut_out11
rlabel metal1 2527 2215 2527 2215 1 lut_out12
rlabel metal1 2998 2214 2998 2214 1 lut_out13
rlabel metal1 3470 2214 3470 2214 1 lut_out14
rlabel metal1 1586 1636 1586 1636 1 lut_out15
rlabel metal1 2057 1636 2057 1636 1 lut_out16
rlabel metal1 2527 1637 2527 1637 1 lut_out17
rlabel metal1 2997 1636 2997 1636 1 lut_out18
rlabel metal1 3469 1636 3469 1636 1 lut_out19
rlabel metal1 1834 3494 1834 3494 1 inp2_1
<< end >>
