magic
tech scmos
timestamp 1414808142
<< nwell >>
rect 16 314 205 371
rect 27 310 54 314
rect 69 310 96 314
<< ntransistor >>
rect 28 276 30 286
rect 36 276 38 296
rect 41 276 43 296
rect 49 276 51 296
rect 54 276 56 296
rect 70 276 72 286
rect 78 276 80 296
rect 83 276 85 296
rect 91 276 93 296
rect 96 276 98 296
rect 112 272 114 292
rect 120 272 122 282
rect 125 272 127 282
rect 134 272 136 282
rect 139 272 141 282
rect 148 272 150 282
rect 164 272 166 282
rect 169 272 171 282
rect 179 272 181 282
rect 184 272 186 282
rect 192 272 194 292
<< ptransistor >>
rect 28 336 30 356
rect 36 316 38 356
rect 41 316 43 356
rect 49 320 51 360
rect 54 320 56 360
rect 70 336 72 356
rect 78 316 80 356
rect 83 316 85 356
rect 91 320 93 360
rect 96 320 98 360
rect 112 320 114 360
rect 120 340 122 360
rect 126 340 128 360
rect 134 340 136 360
rect 140 340 142 360
rect 148 340 150 360
rect 164 340 166 360
rect 169 340 171 360
rect 179 350 181 360
rect 184 350 186 360
rect 192 320 194 360
<< ndiffusion >>
rect 33 294 36 296
rect 27 276 28 286
rect 30 276 31 286
rect 35 276 36 294
rect 38 276 41 296
rect 43 294 49 296
rect 43 276 44 294
rect 48 276 49 294
rect 51 276 54 296
rect 56 276 57 296
rect 75 294 78 296
rect 69 276 70 286
rect 72 276 73 286
rect 77 276 78 294
rect 80 276 83 296
rect 85 294 91 296
rect 85 276 86 294
rect 90 276 91 294
rect 93 276 96 296
rect 98 276 99 296
rect 107 291 112 292
rect 111 272 112 291
rect 114 291 119 292
rect 114 272 115 291
rect 187 291 192 292
rect 119 272 120 282
rect 122 272 125 282
rect 127 281 134 282
rect 127 272 129 281
rect 133 272 134 281
rect 136 272 139 282
rect 141 281 148 282
rect 141 272 142 281
rect 146 272 148 281
rect 150 281 155 282
rect 150 272 151 281
rect 159 281 164 282
rect 163 272 164 281
rect 166 272 169 282
rect 171 281 179 282
rect 171 272 173 281
rect 177 272 179 281
rect 181 272 184 282
rect 186 272 187 282
rect 191 272 192 291
rect 194 291 199 292
rect 194 272 195 291
<< pdiffusion >>
rect 27 336 28 356
rect 30 336 31 356
rect 35 322 36 356
rect 33 316 36 322
rect 38 316 41 356
rect 43 322 44 356
rect 48 322 49 360
rect 43 320 49 322
rect 51 320 54 360
rect 56 320 57 360
rect 69 336 70 356
rect 72 336 73 356
rect 43 316 46 320
rect 77 322 78 356
rect 75 316 78 322
rect 80 316 83 356
rect 85 322 86 356
rect 90 322 91 360
rect 85 320 91 322
rect 93 320 96 360
rect 98 320 99 360
rect 107 359 112 360
rect 111 320 112 359
rect 114 321 115 360
rect 119 340 120 360
rect 122 340 126 360
rect 128 359 134 360
rect 128 340 129 359
rect 133 340 134 359
rect 136 340 140 360
rect 142 359 148 360
rect 142 340 143 359
rect 147 340 148 359
rect 150 359 155 360
rect 150 340 151 359
rect 159 359 164 360
rect 163 340 164 359
rect 166 340 169 360
rect 171 359 179 360
rect 171 340 173 359
rect 177 350 179 359
rect 181 350 184 360
rect 186 359 192 360
rect 186 350 187 359
rect 177 340 178 350
rect 114 320 119 321
rect 85 316 88 320
rect 191 320 192 359
rect 194 359 199 360
rect 194 320 195 359
<< ndcontact >>
rect 23 276 27 286
rect 31 276 35 294
rect 44 276 48 294
rect 57 276 61 296
rect 65 276 69 286
rect 73 276 77 294
rect 86 276 90 294
rect 99 276 103 296
rect 107 272 111 291
rect 115 272 119 291
rect 129 272 133 281
rect 142 272 146 281
rect 151 272 155 281
rect 159 272 163 281
rect 173 272 177 281
rect 187 272 191 291
rect 195 272 199 291
<< pdcontact >>
rect 23 336 27 356
rect 31 322 35 356
rect 44 322 48 360
rect 57 320 61 360
rect 65 336 69 356
rect 73 322 77 356
rect 86 322 90 360
rect 99 320 103 360
rect 107 320 111 359
rect 115 321 119 360
rect 129 340 133 359
rect 143 340 147 359
rect 151 340 155 359
rect 159 340 163 359
rect 173 340 177 359
rect 187 320 191 359
rect 195 320 199 359
<< psubstratepcontact >>
rect 19 264 23 268
rect 35 264 39 268
rect 51 264 55 268
rect 61 264 65 268
rect 77 264 81 268
rect 93 264 97 268
rect 103 264 107 268
rect 119 264 123 268
rect 135 264 139 268
rect 151 264 155 268
rect 167 264 171 268
rect 183 264 187 268
<< nsubstratencontact >>
rect 19 364 23 368
rect 35 364 39 368
rect 51 364 55 368
rect 61 364 65 368
rect 77 364 81 368
rect 93 364 97 368
rect 103 364 107 368
rect 119 364 123 368
rect 135 364 139 368
rect 151 364 155 368
rect 167 364 171 368
rect 183 364 187 368
<< polysilicon >>
rect 28 361 43 363
rect 28 356 30 361
rect 36 356 38 358
rect 41 356 43 361
rect 49 360 51 362
rect 54 360 56 362
rect 70 361 85 363
rect 28 335 30 336
rect 25 333 30 335
rect 25 315 27 333
rect 70 356 72 361
rect 78 356 80 358
rect 83 356 85 361
rect 91 360 93 362
rect 96 360 98 362
rect 112 360 114 362
rect 120 360 122 362
rect 126 360 128 362
rect 134 360 136 362
rect 140 360 142 362
rect 148 360 150 362
rect 164 360 166 362
rect 169 360 171 362
rect 179 360 181 362
rect 184 360 186 362
rect 192 360 194 362
rect 70 335 72 336
rect 67 333 72 335
rect 36 315 38 316
rect 24 313 27 315
rect 32 313 38 315
rect 41 314 43 316
rect 24 309 26 313
rect 32 309 34 313
rect 49 306 51 320
rect 54 319 56 320
rect 54 317 57 319
rect 24 301 26 305
rect 24 299 27 301
rect 25 289 27 299
rect 32 299 34 305
rect 46 304 51 306
rect 41 300 45 302
rect 32 297 38 299
rect 36 296 38 297
rect 41 296 43 300
rect 55 299 57 313
rect 67 309 69 333
rect 78 315 80 316
rect 75 313 80 315
rect 83 314 85 316
rect 75 309 77 313
rect 91 306 93 320
rect 96 319 98 320
rect 96 317 99 319
rect 49 296 51 298
rect 54 297 57 299
rect 54 296 56 297
rect 25 287 30 289
rect 28 286 30 287
rect 67 289 69 305
rect 74 299 76 305
rect 88 304 93 306
rect 83 300 87 302
rect 74 297 80 299
rect 78 296 80 297
rect 83 296 85 300
rect 97 299 99 313
rect 112 303 114 320
rect 120 312 122 340
rect 91 296 93 298
rect 96 297 99 299
rect 96 296 98 297
rect 67 287 72 289
rect 70 286 72 287
rect 112 292 114 299
rect 28 271 30 276
rect 36 274 38 276
rect 41 274 43 276
rect 49 271 51 276
rect 54 274 56 276
rect 28 269 51 271
rect 70 271 72 276
rect 78 274 80 276
rect 83 274 85 276
rect 91 271 93 276
rect 96 274 98 276
rect 120 282 122 308
rect 126 304 128 340
rect 134 320 136 340
rect 134 295 136 316
rect 125 293 136 295
rect 140 337 142 340
rect 125 282 127 293
rect 140 289 142 333
rect 148 327 150 340
rect 164 339 166 340
rect 155 337 166 339
rect 135 285 136 289
rect 134 282 136 285
rect 139 285 140 289
rect 139 282 141 285
rect 148 282 150 323
rect 154 285 156 333
rect 169 329 171 340
rect 179 333 181 350
rect 177 331 181 333
rect 164 327 171 329
rect 162 290 164 299
rect 169 297 171 327
rect 184 319 186 350
rect 180 317 186 319
rect 179 297 181 313
rect 192 311 194 320
rect 190 307 194 311
rect 169 295 176 297
rect 162 288 171 290
rect 154 283 166 285
rect 164 282 166 283
rect 169 282 171 288
rect 174 285 176 295
rect 179 293 180 297
rect 174 283 181 285
rect 179 282 181 283
rect 184 282 186 297
rect 192 292 194 307
rect 70 269 93 271
rect 112 270 114 272
rect 120 270 122 272
rect 125 270 127 272
rect 134 270 136 272
rect 139 270 141 272
rect 148 270 150 272
rect 164 270 166 272
rect 169 270 171 272
rect 179 270 181 272
rect 184 270 186 272
rect 192 270 194 272
<< polycontact >>
rect 22 305 26 309
rect 30 305 34 309
rect 42 302 46 306
rect 55 313 59 317
rect 65 305 69 309
rect 73 305 77 309
rect 84 302 88 306
rect 97 313 101 317
rect 118 308 122 312
rect 111 299 115 303
rect 132 316 136 320
rect 126 300 130 304
rect 140 333 144 337
rect 146 323 150 327
rect 131 285 135 289
rect 140 285 144 289
rect 154 333 158 337
rect 160 325 164 329
rect 175 327 179 331
rect 160 299 164 303
rect 178 313 182 317
rect 186 307 190 311
rect 180 293 184 297
<< metal1 >>
rect 34 372 195 376
rect 19 368 203 369
rect 23 364 35 368
rect 39 364 51 368
rect 55 364 61 368
rect 65 364 77 368
rect 81 364 93 368
rect 97 364 103 368
rect 107 364 119 368
rect 123 364 135 368
rect 139 364 151 368
rect 155 364 167 368
rect 171 364 183 368
rect 187 364 203 368
rect 19 363 203 364
rect 31 356 35 363
rect 57 360 61 363
rect 23 319 26 336
rect 48 322 52 325
rect 23 316 42 319
rect 22 309 26 313
rect 39 302 42 316
rect 49 303 52 322
rect 73 356 77 363
rect 99 360 103 363
rect 115 360 119 363
rect 65 319 68 336
rect 90 322 94 325
rect 65 316 84 319
rect 65 309 69 313
rect 39 300 44 302
rect 23 297 44 300
rect 49 299 58 303
rect 81 302 84 316
rect 91 303 94 322
rect 107 359 111 360
rect 103 320 104 323
rect 100 317 104 320
rect 101 313 104 317
rect 129 359 133 360
rect 123 340 129 343
rect 143 359 147 363
rect 151 359 155 360
rect 159 359 163 363
rect 172 359 178 360
rect 172 340 173 359
rect 177 340 178 359
rect 187 359 191 363
rect 151 337 154 340
rect 144 334 154 337
rect 127 323 146 326
rect 153 326 160 329
rect 153 320 156 326
rect 172 322 175 331
rect 111 316 132 318
rect 136 317 156 320
rect 163 319 175 322
rect 195 359 199 360
rect 107 315 135 316
rect 115 310 118 312
rect 104 307 118 310
rect 104 303 107 307
rect 81 300 86 302
rect 23 286 26 297
rect 49 296 52 299
rect 67 297 86 300
rect 91 299 107 303
rect 115 300 126 303
rect 163 303 166 319
rect 195 317 199 320
rect 182 314 195 317
rect 175 307 186 310
rect 130 300 160 303
rect 48 291 52 296
rect 67 290 70 297
rect 91 296 94 299
rect 66 286 70 290
rect 90 291 94 296
rect 31 269 35 276
rect 57 269 61 276
rect 73 269 77 276
rect 99 269 103 276
rect 107 291 111 292
rect 115 291 119 292
rect 132 289 135 300
rect 164 300 166 303
rect 195 297 199 313
rect 184 294 199 297
rect 195 291 199 294
rect 144 285 154 288
rect 151 282 154 285
rect 123 281 133 282
rect 123 279 129 281
rect 142 281 147 282
rect 146 272 147 281
rect 151 281 155 282
rect 159 281 163 282
rect 171 281 178 282
rect 171 279 173 281
rect 172 272 173 279
rect 177 272 178 281
rect 115 269 119 272
rect 142 269 147 272
rect 159 269 163 272
rect 187 269 191 272
rect 19 268 203 269
rect 23 264 35 268
rect 39 264 51 268
rect 55 264 61 268
rect 65 264 77 268
rect 81 264 93 268
rect 97 264 103 268
rect 107 264 119 268
rect 123 264 135 268
rect 139 264 151 268
rect 155 264 167 268
rect 171 264 183 268
rect 187 264 203 268
rect 19 263 203 264
rect 62 256 73 260
<< m2contact >>
rect 30 372 34 376
rect 195 372 199 376
rect 30 309 34 313
rect 73 309 77 313
rect 58 299 62 303
rect 123 336 127 340
rect 171 336 175 340
rect 123 323 127 327
rect 107 316 111 320
rect 195 313 199 317
rect 171 306 175 310
rect 107 292 111 296
rect 123 282 127 286
rect 171 282 175 286
rect 58 256 62 260
rect 73 256 77 260
<< metal2 >>
rect 30 313 34 372
rect 123 327 127 336
rect 58 260 62 299
rect 73 260 77 309
rect 107 296 111 316
rect 123 286 127 323
rect 171 310 175 336
rect 195 317 199 372
rect 171 286 175 306
<< m1p >>
rect 22 309 26 313
rect 30 309 34 313
rect 55 309 59 313
rect 65 309 69 313
rect 195 309 199 313
rect 115 299 119 303
<< labels >>
rlabel metal1 117 300 117 300 1 Clk
rlabel metal1 197 310 197 310 1 Q
rlabel metal1 94 300 94 300 1 muxout2
rlabel metal1 25 365 25 365 1 Vdd
rlabel metal1 25 265 25 265 1 Gnd
rlabel metal1 51 300 51 300 1 muxout1
rlabel metal1 67 310 67 310 1 Reset
rlabel polysilicon 57 310 57 310 1 D
rlabel metal1 24 310 24 310 1 Load
<< end >>
