magic
tech scmos
timestamp 1415084864
<< metal1 >>
rect 2342 3992 2354 4004
rect 1008 3980 1334 3992
rect 1346 3980 1805 3992
rect 1817 3980 1910 3992
rect 1922 3980 2276 3992
rect 2288 3980 2743 3992
rect 2755 3980 2809 3992
rect 2821 3980 3218 3992
rect 3230 3980 3992 3992
rect 1008 1020 1020 3980
rect 1028 3960 1043 3972
rect 1055 3960 2156 3972
rect 2168 3960 2542 3972
rect 2554 3960 3055 3972
rect 3067 3960 3143 3972
rect 3155 3960 3972 3972
rect 1028 3651 1040 3960
rect 1872 3761 1946 3765
rect 2656 3761 2761 3765
rect 2814 3761 2846 3765
rect 3127 3761 3359 3765
rect 1250 3754 1818 3758
rect 1822 3754 2269 3758
rect 2273 3754 2659 3758
rect 2663 3754 2760 3758
rect 2764 3754 3130 3758
rect 3134 3754 3343 3758
rect 1326 3745 1334 3751
rect 1813 3745 1820 3751
rect 2739 3745 2747 3751
rect 2755 3745 2766 3751
rect 1318 3714 1363 3718
rect 3202 3714 3248 3718
rect 1851 3681 1864 3685
rect 2793 3681 2806 3685
rect 1239 3671 1250 3675
rect 1327 3669 1378 3673
rect 1860 3671 1864 3681
rect 2802 3671 2806 3681
rect 3215 3669 3262 3673
rect 2735 3666 2740 3667
rect 1048 3659 1227 3664
rect 2324 3661 2652 3665
rect 2735 3664 2736 3666
rect 1882 3654 2209 3658
rect 2309 3654 2652 3658
rect 2824 3654 3097 3658
rect 1028 3645 1248 3651
rect 1326 3645 1814 3651
rect 1876 3645 2661 3651
rect 2739 3645 2770 3651
rect 2818 3645 3216 3651
rect 1028 3453 1040 3645
rect 1328 3638 1350 3642
rect 1763 3638 1821 3642
rect 2234 3638 2293 3642
rect 2705 3638 2764 3642
rect 3176 3638 3234 3642
rect 1327 3629 1334 3635
rect 3101 3624 3151 3628
rect 1232 3593 1242 3597
rect 1263 3575 1267 3593
rect 1239 3559 1247 3563
rect 1326 3514 1332 3535
rect 1326 3508 1346 3514
rect 1324 3493 1345 3497
rect 1742 3493 1816 3497
rect 2684 3493 2758 3497
rect 1028 1040 1040 3441
rect 1241 3362 1354 3366
rect 2213 3362 2287 3366
rect 3155 3362 3229 3366
rect 3626 3239 3702 3243
rect 1317 3102 1350 3106
rect 1763 3102 1821 3106
rect 2234 3102 2292 3106
rect 2705 3102 2763 3106
rect 3176 3102 3233 3106
rect 3644 3088 3772 3092
rect 1275 3081 1355 3085
rect 1366 3081 1738 3085
rect 1836 3081 2209 3085
rect 2310 3081 2680 3085
rect 2779 3081 3151 3085
rect 3252 3081 3622 3085
rect 1275 3074 1738 3078
rect 1838 3074 2680 3078
rect 2781 3074 3622 3078
rect 1382 3067 1518 3071
rect 1614 3067 1875 3071
rect 1889 3067 1977 3071
rect 2085 3067 2299 3071
rect 2324 3067 2460 3071
rect 2556 3067 2819 3071
rect 2831 3067 2919 3071
rect 3027 3067 3239 3071
rect 3266 3067 3402 3071
rect 1621 3060 1764 3064
rect 2093 3060 2235 3064
rect 2564 3060 2706 3064
rect 3034 3060 3177 3064
rect 3494 3060 3597 3064
rect 3566 3046 3643 3050
rect 1764 2517 1788 2521
rect 2235 2517 2259 2521
rect 2706 2517 2730 2521
rect 3177 2517 3201 2521
rect 3647 2517 3746 2521
rect 1784 2510 1788 2517
rect 2255 2510 2259 2517
rect 2726 2510 2730 2517
rect 3197 2510 3201 2517
rect 1366 2503 2209 2507
rect 2308 2503 3151 2507
rect 3250 2503 3747 2507
rect 1366 2496 1738 2500
rect 1837 2496 2209 2500
rect 2310 2496 2680 2500
rect 2779 2496 3151 2500
rect 3252 2496 3622 2500
rect 1382 2489 1518 2493
rect 1889 2489 1977 2493
rect 2324 2489 2460 2493
rect 2831 2489 2919 2493
rect 3266 2489 3402 2493
rect 1245 2482 1354 2486
rect 1763 2482 1821 2486
rect 2234 2482 2300 2486
rect 2705 2482 2774 2486
rect 3176 2482 3234 2486
rect 1742 2337 1816 2341
rect 2684 2337 2758 2341
rect 1245 2206 1356 2210
rect 2213 2206 2287 2210
rect 3155 2206 3229 2210
rect 3642 2003 3765 2007
rect 1317 1946 1350 1950
rect 1763 1946 1821 1950
rect 2234 1946 2291 1950
rect 2705 1946 2763 1950
rect 3176 1946 3234 1950
rect 3643 1932 3758 1936
rect 1366 1925 1738 1929
rect 1837 1925 2209 1929
rect 2309 1925 2680 1929
rect 2779 1925 3151 1929
rect 3252 1925 3622 1929
rect 1233 1918 1738 1922
rect 1839 1918 2680 1922
rect 2781 1918 3622 1922
rect 1233 1911 1355 1915
rect 1382 1911 1518 1915
rect 1614 1911 1878 1915
rect 1889 1911 1977 1915
rect 2085 1911 2297 1915
rect 2324 1911 2460 1915
rect 2556 1911 2820 1915
rect 2831 1911 2919 1915
rect 3027 1911 3241 1915
rect 3266 1911 3402 1915
rect 1621 1904 1764 1908
rect 2093 1904 2235 1908
rect 2563 1904 2706 1908
rect 3035 1904 3177 1908
rect 3494 1904 3597 1908
rect 3565 1890 3643 1894
rect 1764 1361 1784 1365
rect 2235 1361 2255 1365
rect 2705 1361 2726 1365
rect 3177 1361 3201 1365
rect 3647 1361 3729 1365
rect 1317 1354 1319 1358
rect 3197 1354 3201 1361
rect 1366 1347 2209 1351
rect 2308 1347 3151 1351
rect 3250 1347 3730 1351
rect 1658 1340 1738 1344
rect 1837 1340 1890 1344
rect 2622 1340 2680 1344
rect 2779 1340 2830 1344
rect 3503 1340 3622 1344
rect 3960 1040 3972 3960
rect 1028 1028 1766 1040
rect 1778 1028 2237 1040
rect 2249 1028 2642 1040
rect 2654 1028 2708 1040
rect 2720 1028 3179 1040
rect 3191 1028 3650 1040
rect 3662 1028 3972 1040
rect 3980 1020 3992 3980
rect 1008 1008 3992 1020
<< m2contact >>
rect 1334 3980 1346 3992
rect 1805 3980 1817 3992
rect 1910 3980 1922 3992
rect 2276 3980 2288 3992
rect 2743 3980 2755 3992
rect 2809 3980 2821 3992
rect 3218 3980 3230 3992
rect 1043 3960 1055 3972
rect 2156 3960 2168 3972
rect 2542 3960 2554 3972
rect 3055 3960 3067 3972
rect 3143 3960 3155 3972
rect 1868 3761 1872 3765
rect 1946 3761 1951 3766
rect 2652 3761 2656 3765
rect 2761 3761 2766 3766
rect 2810 3761 2814 3765
rect 2846 3761 2851 3766
rect 3123 3761 3127 3765
rect 3359 3761 3364 3766
rect 1246 3754 1250 3758
rect 1818 3754 1822 3758
rect 2269 3754 2273 3758
rect 2659 3754 2663 3758
rect 2760 3754 2764 3758
rect 3130 3754 3134 3758
rect 1334 3743 1342 3751
rect 1805 3743 1813 3751
rect 2276 3743 2284 3751
rect 2747 3743 2755 3751
rect 1363 3714 1367 3718
rect 1868 3715 1872 3719
rect 2810 3713 2814 3717
rect 3248 3714 3252 3718
rect 1826 3691 1830 3695
rect 1850 3691 1854 3695
rect 2269 3691 2273 3695
rect 2768 3691 2772 3695
rect 2792 3691 2796 3695
rect 1235 3671 1239 3675
rect 1378 3669 1382 3673
rect 3211 3669 3215 3673
rect 3262 3669 3266 3673
rect 1043 3659 1048 3664
rect 1227 3659 1232 3664
rect 2320 3661 2324 3665
rect 2652 3661 2656 3665
rect 2736 3662 2740 3666
rect 1878 3654 1882 3658
rect 2209 3654 2213 3658
rect 2305 3654 2309 3658
rect 2652 3654 2656 3658
rect 2820 3654 2824 3658
rect 3097 3654 3101 3658
rect 1324 3638 1328 3642
rect 1334 3627 1342 3635
rect 1777 3631 1781 3635
rect 2248 3631 2252 3635
rect 2719 3631 2723 3635
rect 3190 3631 3194 3635
rect 3661 3631 3665 3635
rect 3097 3624 3101 3628
rect 3151 3624 3155 3628
rect 1227 3592 1232 3597
rect 1242 3593 1246 3597
rect 1263 3593 1267 3597
rect 1235 3559 1239 3563
rect 1320 3546 1324 3550
rect 1784 3501 1788 3505
rect 2255 3501 2259 3505
rect 2726 3501 2730 3505
rect 3197 3501 3201 3505
rect 3668 3501 3672 3505
rect 1320 3493 1324 3497
rect 1363 3493 1367 3497
rect 1738 3493 1742 3497
rect 2305 3493 2309 3497
rect 2680 3493 2684 3497
rect 3248 3493 3252 3497
rect 1028 3441 1040 3453
rect 2209 3362 2213 3366
rect 2775 3362 2779 3366
rect 3151 3362 3155 3366
rect 3622 3239 3626 3243
rect 1738 3181 1742 3185
rect 2209 3181 2213 3185
rect 2680 3181 2684 3185
rect 3151 3181 3155 3185
rect 3622 3181 3626 3185
rect 1738 3151 1742 3155
rect 2680 3151 2684 3155
rect 3622 3151 3626 3155
rect 1327 3116 1331 3120
rect 1798 3116 1802 3120
rect 2269 3116 2273 3120
rect 2740 3116 2744 3120
rect 3211 3116 3215 3120
rect 1313 3102 1317 3106
rect 1759 3102 1763 3106
rect 2230 3102 2234 3106
rect 2701 3102 2705 3106
rect 3172 3102 3176 3106
rect 1320 3095 1324 3099
rect 1791 3095 1795 3099
rect 2262 3095 2266 3099
rect 2733 3095 2737 3099
rect 3204 3095 3208 3099
rect 1758 3088 1762 3092
rect 2230 3088 2234 3092
rect 2701 3088 2705 3092
rect 3172 3088 3176 3092
rect 1355 3081 1359 3085
rect 1362 3081 1366 3085
rect 1738 3081 1742 3085
rect 1832 3081 1836 3085
rect 2209 3081 2213 3085
rect 2306 3081 2310 3085
rect 2680 3081 2684 3085
rect 2775 3081 2779 3085
rect 3151 3081 3155 3085
rect 3248 3081 3252 3085
rect 3622 3081 3626 3085
rect 1738 3074 1742 3078
rect 1834 3074 1838 3078
rect 2680 3074 2684 3078
rect 2777 3074 2781 3078
rect 3622 3074 3626 3078
rect 1378 3067 1382 3071
rect 1518 3067 1522 3071
rect 1610 3067 1614 3071
rect 1875 3067 1879 3071
rect 1885 3067 1889 3071
rect 1977 3067 1981 3071
rect 2081 3067 2085 3071
rect 2299 3067 2303 3071
rect 2320 3067 2324 3071
rect 2460 3067 2464 3071
rect 2552 3067 2556 3071
rect 2819 3067 2823 3071
rect 2827 3067 2831 3071
rect 2919 3067 2923 3071
rect 3023 3067 3027 3071
rect 3239 3067 3243 3071
rect 3262 3067 3266 3071
rect 3402 3067 3406 3071
rect 1617 3060 1621 3064
rect 2089 3060 2093 3064
rect 2560 3060 2564 3064
rect 3030 3060 3034 3064
rect 3597 3060 3601 3064
rect 1777 3053 1781 3057
rect 2248 3053 2252 3057
rect 2719 3053 2723 3057
rect 3190 3053 3194 3057
rect 3661 3053 3665 3057
rect 3562 3046 3566 3050
rect 3643 3046 3647 3050
rect 1784 2923 1788 2927
rect 2255 2923 2259 2927
rect 2726 2923 2730 2927
rect 3197 2923 3201 2927
rect 3668 2923 3672 2927
rect 1362 2915 1366 2919
rect 1834 2915 1838 2919
rect 2306 2915 2310 2919
rect 2777 2915 2781 2919
rect 3248 2915 3252 2919
rect 1362 2784 1366 2788
rect 1833 2784 1837 2788
rect 2304 2784 2308 2788
rect 2775 2784 2779 2788
rect 3246 2784 3250 2788
rect 1738 2603 1742 2607
rect 2209 2603 2213 2607
rect 2680 2603 2684 2607
rect 3151 2603 3155 2607
rect 3622 2603 3626 2607
rect 1738 2573 1742 2577
rect 2209 2573 2213 2577
rect 2680 2573 2684 2577
rect 3151 2573 3155 2577
rect 3622 2573 3626 2577
rect 1327 2538 1331 2542
rect 1798 2538 1802 2542
rect 2269 2538 2273 2542
rect 2740 2538 2744 2542
rect 3211 2538 3215 2542
rect 1320 2517 1324 2521
rect 1791 2517 1795 2521
rect 2262 2517 2266 2521
rect 2733 2517 2737 2521
rect 3204 2517 3208 2521
rect 1313 2510 1317 2514
rect 1362 2503 1366 2507
rect 2209 2503 2213 2507
rect 2304 2503 2308 2507
rect 3151 2503 3155 2507
rect 3246 2503 3250 2507
rect 1362 2496 1366 2500
rect 1738 2496 1742 2500
rect 1833 2496 1837 2500
rect 2209 2496 2213 2500
rect 2306 2496 2310 2500
rect 2680 2496 2684 2500
rect 2775 2496 2779 2500
rect 3151 2496 3155 2500
rect 3248 2496 3252 2500
rect 3622 2496 3626 2500
rect 1378 2489 1382 2493
rect 1518 2489 1522 2493
rect 1885 2489 1889 2493
rect 1977 2489 1981 2493
rect 2320 2489 2324 2493
rect 2460 2489 2464 2493
rect 2827 2489 2831 2493
rect 2919 2489 2923 2493
rect 3262 2489 3266 2493
rect 3402 2489 3406 2493
rect 1777 2475 1781 2479
rect 2248 2475 2252 2479
rect 2719 2475 2723 2479
rect 3190 2475 3194 2479
rect 3661 2475 3665 2479
rect 1784 2345 1788 2349
rect 2255 2345 2259 2349
rect 2726 2345 2730 2349
rect 3197 2345 3201 2349
rect 3668 2345 3672 2349
rect 1362 2337 1366 2341
rect 1738 2337 1742 2341
rect 2306 2337 2310 2341
rect 2680 2337 2684 2341
rect 3248 2337 3252 2341
rect 1833 2206 1837 2210
rect 2209 2206 2213 2210
rect 2775 2206 2779 2210
rect 3151 2206 3155 2210
rect 1738 2025 1742 2029
rect 2209 2025 2213 2029
rect 2680 2025 2684 2029
rect 3151 2025 3155 2029
rect 1738 1995 1742 1999
rect 2680 1995 2684 1999
rect 3622 1995 3626 1999
rect 1327 1960 1331 1964
rect 1798 1960 1802 1964
rect 2269 1960 2273 1964
rect 2740 1960 2744 1964
rect 3211 1960 3215 1964
rect 1313 1946 1317 1950
rect 1759 1946 1763 1950
rect 2230 1946 2234 1950
rect 2701 1946 2705 1950
rect 3172 1946 3176 1950
rect 1320 1939 1324 1943
rect 1791 1939 1795 1943
rect 2262 1939 2266 1943
rect 2733 1939 2737 1943
rect 3204 1939 3208 1943
rect 1759 1932 1763 1936
rect 2230 1932 2234 1936
rect 2701 1932 2705 1936
rect 3172 1932 3176 1936
rect 1362 1925 1366 1929
rect 1738 1925 1742 1929
rect 1833 1925 1837 1929
rect 2209 1925 2213 1929
rect 2305 1925 2309 1929
rect 2680 1925 2684 1929
rect 2775 1925 2779 1929
rect 3151 1925 3155 1929
rect 3248 1925 3252 1929
rect 3622 1925 3626 1929
rect 1738 1918 1742 1922
rect 1835 1918 1839 1922
rect 2680 1918 2684 1922
rect 2777 1918 2781 1922
rect 3622 1918 3626 1922
rect 1355 1911 1359 1915
rect 1378 1911 1382 1915
rect 1518 1911 1522 1915
rect 1610 1911 1614 1915
rect 1878 1911 1882 1915
rect 1885 1911 1889 1915
rect 1977 1911 1981 1915
rect 2081 1911 2085 1915
rect 2297 1911 2301 1915
rect 2320 1911 2324 1915
rect 2460 1911 2464 1915
rect 2552 1911 2556 1915
rect 2820 1911 2824 1915
rect 2827 1911 2831 1915
rect 2919 1911 2923 1915
rect 3023 1911 3027 1915
rect 3241 1911 3245 1915
rect 3262 1911 3266 1915
rect 3402 1911 3406 1915
rect 1617 1904 1621 1908
rect 2089 1904 2093 1908
rect 2559 1904 2563 1908
rect 3031 1904 3035 1908
rect 3597 1904 3601 1908
rect 1777 1897 1781 1901
rect 2248 1897 2252 1901
rect 2719 1897 2723 1901
rect 3190 1897 3194 1901
rect 3661 1897 3665 1901
rect 3561 1890 3565 1894
rect 3643 1890 3647 1894
rect 1784 1767 1788 1771
rect 2255 1767 2259 1771
rect 2726 1767 2730 1771
rect 3197 1767 3201 1771
rect 3668 1767 3672 1771
rect 1362 1759 1366 1763
rect 1835 1759 1839 1763
rect 2305 1759 2309 1763
rect 2777 1759 2781 1763
rect 3248 1759 3252 1763
rect 1362 1628 1366 1632
rect 1833 1628 1837 1632
rect 2304 1628 2308 1632
rect 2775 1628 2779 1632
rect 3246 1628 3250 1632
rect 1738 1447 1742 1451
rect 2209 1447 2213 1451
rect 2680 1447 2684 1451
rect 3151 1447 3155 1451
rect 3622 1447 3626 1451
rect 1738 1417 1742 1421
rect 2209 1417 2213 1421
rect 2680 1417 2684 1421
rect 3151 1417 3155 1421
rect 3622 1417 3626 1421
rect 1327 1382 1331 1386
rect 1798 1382 1802 1386
rect 2269 1382 2273 1386
rect 2740 1382 2744 1386
rect 3211 1382 3215 1386
rect 1320 1361 1324 1365
rect 1784 1361 1788 1365
rect 1791 1361 1795 1365
rect 2255 1361 2259 1365
rect 2262 1361 2266 1365
rect 2726 1361 2730 1365
rect 2733 1361 2737 1365
rect 3204 1361 3208 1365
rect 1313 1354 1317 1358
rect 1784 1354 1788 1358
rect 2255 1354 2259 1358
rect 2726 1354 2730 1358
rect 1362 1347 1366 1351
rect 2209 1347 2213 1351
rect 2304 1347 2308 1351
rect 3151 1347 3155 1351
rect 3246 1347 3250 1351
rect 1654 1340 1658 1344
rect 1738 1340 1742 1344
rect 1833 1340 1837 1344
rect 1890 1340 1894 1344
rect 2618 1340 2622 1344
rect 2680 1340 2684 1344
rect 2775 1340 2779 1344
rect 2830 1340 2834 1344
rect 3499 1340 3503 1344
rect 3622 1340 3626 1344
rect 1766 1028 1778 1040
rect 2237 1028 2249 1040
rect 2642 1028 2654 1040
rect 2708 1028 2720 1040
rect 3179 1028 3191 1040
rect 3650 1028 3662 1040
<< metal2 >>
rect 1011 3995 1020 4000
rect 1044 3995 1053 4000
rect 1011 3986 1053 3995
rect 1044 3972 1053 3986
rect 1259 3770 1264 4000
rect 1911 3992 1920 4000
rect 1236 3765 1264 3770
rect 1236 3695 1241 3765
rect 1246 3706 1250 3754
rect 1334 3751 1342 3980
rect 1000 3659 1043 3664
rect 1227 3597 1232 3659
rect 1235 3563 1239 3671
rect 1322 3669 1331 3673
rect 1246 3593 1263 3597
rect 1242 3579 1246 3583
rect 1324 3553 1328 3638
rect 1334 3635 1342 3743
rect 1805 3751 1813 3980
rect 1946 3766 1951 4009
rect 2157 3972 2166 4000
rect 2511 3995 2520 4000
rect 2544 3995 2553 4000
rect 2511 3986 2553 3995
rect 1320 3497 1324 3546
rect 1000 3444 1028 3453
rect 1005 3420 1014 3444
rect 1000 3411 1014 3420
rect 1313 2514 1317 3102
rect 1320 2521 1324 3095
rect 1313 1358 1317 1946
rect 1320 1943 1324 2517
rect 1320 1365 1324 1939
rect 1327 2542 1331 3116
rect 1327 1964 1331 2538
rect 1327 1386 1331 1960
rect 1334 1496 1342 3627
rect 1363 3497 1367 3714
rect 1378 3638 1382 3669
rect 1738 3185 1742 3493
rect 1355 3092 1425 3096
rect 1355 3085 1359 3092
rect 1362 2919 1366 3081
rect 1421 3060 1425 3092
rect 1738 3085 1742 3151
rect 1759 3092 1763 3102
rect 1762 3088 1763 3092
rect 1525 3078 1621 3082
rect 1525 3060 1529 3078
rect 1610 3060 1614 3067
rect 1617 3064 1621 3078
rect 1421 3056 1529 3060
rect 1362 2507 1366 2784
rect 1738 2607 1742 3074
rect 1738 2500 1742 2573
rect 1362 2341 1366 2496
rect 1738 2029 1742 2337
rect 1355 1936 1425 1940
rect 1355 1915 1359 1936
rect 1362 1763 1366 1925
rect 1421 1904 1425 1936
rect 1738 1929 1742 1995
rect 1759 1936 1763 1946
rect 1525 1922 1621 1926
rect 1525 1904 1529 1922
rect 1610 1904 1614 1911
rect 1617 1908 1621 1922
rect 1421 1900 1529 1904
rect 1362 1351 1366 1628
rect 1738 1451 1742 1918
rect 1738 1344 1742 1417
rect 1518 1293 1522 1339
rect 1654 1293 1658 1340
rect 1766 1040 1774 3508
rect 1777 3057 1781 3631
rect 1777 2479 1781 3053
rect 1777 1901 1781 2475
rect 1784 2927 1788 3501
rect 1784 2349 1788 2923
rect 1784 1771 1788 2345
rect 1791 2521 1795 3095
rect 1791 1943 1795 2517
rect 1791 1365 1795 1939
rect 1798 2542 1802 3116
rect 1798 1964 1802 2538
rect 1798 1386 1802 1960
rect 1805 1496 1813 3743
rect 1818 3691 1822 3754
rect 1868 3719 1872 3761
rect 2269 3695 2273 3754
rect 1854 3691 1889 3695
rect 2276 3751 2284 3980
rect 2544 3972 2553 3986
rect 1826 3658 1830 3691
rect 1826 3654 1878 3658
rect 1885 3629 1889 3691
rect 2209 3366 2213 3654
rect 1832 3085 1836 3366
rect 2209 3185 2213 3362
rect 2230 3092 2234 3102
rect 1875 3078 1897 3082
rect 1834 2919 1838 3074
rect 1875 3071 1879 3078
rect 1885 3062 1889 3067
rect 1893 3060 1897 3078
rect 1998 3078 2093 3082
rect 1998 3060 2002 3078
rect 2081 3060 2085 3067
rect 2089 3064 2093 3078
rect 1893 3056 2002 3060
rect 1833 2500 1837 2784
rect 2209 2607 2213 3081
rect 2209 2507 2213 2573
rect 1885 2482 1889 2489
rect 2209 2210 2213 2496
rect 1833 1929 1837 2206
rect 2209 2029 2213 2206
rect 2230 1936 2234 1946
rect 1878 1922 1896 1926
rect 1835 1763 1839 1918
rect 1878 1915 1882 1922
rect 1885 1905 1889 1911
rect 1892 1904 1896 1922
rect 1997 1922 2093 1926
rect 1997 1904 2001 1922
rect 2081 1904 2085 1911
rect 2089 1908 2093 1922
rect 1892 1900 2001 1904
rect 1784 1358 1788 1361
rect 1833 1344 1837 1628
rect 2209 1451 2213 1925
rect 2209 1351 2213 1417
rect 1890 1283 1894 1340
rect 1977 1283 1981 1341
rect 2237 1040 2245 3508
rect 2248 3057 2252 3631
rect 2248 2479 2252 3053
rect 2248 1901 2252 2475
rect 2255 2927 2259 3501
rect 2255 2349 2259 2923
rect 2255 1771 2259 2345
rect 2262 2521 2266 3095
rect 2262 1943 2266 2517
rect 2262 1365 2266 1939
rect 2269 2542 2273 3116
rect 2269 1964 2273 2538
rect 2269 1386 2273 1960
rect 2276 1495 2284 3743
rect 2652 3695 2656 3761
rect 2659 3706 2663 3754
rect 2747 3751 2755 3980
rect 2761 3766 2766 4009
rect 2811 3992 2820 4000
rect 2846 3766 2851 4000
rect 3057 3972 3066 4000
rect 3111 3994 3120 4000
rect 3144 3994 3153 4000
rect 3111 3985 3153 3994
rect 3144 3972 3153 3985
rect 2652 3669 2704 3673
rect 2652 3665 2656 3669
rect 2305 3497 2309 3654
rect 2320 3636 2324 3661
rect 2736 3658 2740 3662
rect 2656 3654 2740 3658
rect 2680 3185 2684 3493
rect 2299 3092 2372 3096
rect 2299 3071 2303 3092
rect 2306 2919 2310 3081
rect 2368 3060 2372 3092
rect 2680 3085 2684 3151
rect 2701 3092 2705 3102
rect 2468 3078 2564 3082
rect 2468 3060 2472 3078
rect 2552 3060 2556 3067
rect 2560 3064 2564 3078
rect 2368 3056 2472 3060
rect 2304 2507 2308 2784
rect 2680 2607 2684 3074
rect 2680 2500 2684 2573
rect 2306 2341 2310 2496
rect 2680 2029 2684 2337
rect 2297 1936 2367 1940
rect 2297 1915 2301 1936
rect 2305 1763 2309 1925
rect 2363 1904 2367 1936
rect 2680 1929 2684 1995
rect 2701 1936 2705 1946
rect 2467 1922 2563 1926
rect 2467 1904 2471 1922
rect 2552 1904 2556 1911
rect 2559 1908 2563 1922
rect 2363 1900 2471 1904
rect 2255 1358 2259 1361
rect 2304 1351 2308 1628
rect 2680 1451 2684 1918
rect 2680 1344 2684 1417
rect 2460 1280 2464 1337
rect 2618 1280 2622 1340
rect 2708 1040 2716 3508
rect 2719 3057 2723 3631
rect 2719 2479 2723 3053
rect 2719 1901 2723 2475
rect 2726 2927 2730 3501
rect 2726 2349 2730 2923
rect 2726 1771 2730 2345
rect 2733 2521 2737 3095
rect 2733 1943 2737 2517
rect 2733 1365 2737 1939
rect 2740 2542 2744 3116
rect 2740 1964 2744 2538
rect 2740 1386 2744 1960
rect 2747 1495 2755 3743
rect 2760 3691 2764 3754
rect 2810 3717 2814 3761
rect 3123 3695 3127 3761
rect 3130 3706 3134 3754
rect 2796 3691 2831 3695
rect 2768 3658 2772 3691
rect 2768 3654 2820 3658
rect 2827 3638 2831 3691
rect 3207 3669 3211 3673
rect 3097 3628 3101 3654
rect 3151 3366 3155 3624
rect 2775 3085 2779 3362
rect 3151 3185 3155 3362
rect 3172 3092 3176 3102
rect 2819 3078 2843 3082
rect 2777 2919 2781 3074
rect 2819 3071 2823 3078
rect 2827 3060 2831 3067
rect 2839 3061 2843 3078
rect 2942 3078 3034 3082
rect 2942 3061 2946 3078
rect 2839 3057 2946 3061
rect 3023 3060 3027 3067
rect 3030 3064 3034 3078
rect 2775 2500 2779 2784
rect 3151 2607 3155 3081
rect 3151 2507 3155 2573
rect 2827 2482 2831 2489
rect 3151 2210 3155 2496
rect 2775 1929 2779 2206
rect 3151 2029 3155 2206
rect 3172 1936 3176 1946
rect 2820 1922 2838 1926
rect 2777 1763 2781 1918
rect 2820 1915 2824 1922
rect 2827 1898 2831 1911
rect 2834 1904 2838 1922
rect 2938 1922 3035 1926
rect 2938 1904 2942 1922
rect 3023 1904 3027 1911
rect 3031 1908 3035 1922
rect 2834 1900 2942 1904
rect 2726 1358 2730 1361
rect 2775 1344 2779 1628
rect 3151 1451 3155 1925
rect 3151 1351 3155 1417
rect 2830 1292 2834 1340
rect 2919 1292 2923 1338
rect 3179 1040 3187 3273
rect 3190 3057 3194 3631
rect 3190 2479 3194 3053
rect 3190 1901 3194 2475
rect 3197 2927 3201 3501
rect 3197 2349 3201 2923
rect 3197 1771 3201 2345
rect 3204 2521 3208 3095
rect 3204 1943 3208 2517
rect 3204 1365 3208 1939
rect 3211 2542 3215 3116
rect 3211 1964 3215 2538
rect 3211 1386 3215 1960
rect 3218 1495 3226 3980
rect 3359 3766 3364 4000
rect 3248 3497 3252 3714
rect 3262 3645 3266 3669
rect 3622 3185 3626 3239
rect 3239 3091 3315 3095
rect 3239 3071 3243 3091
rect 3248 2919 3252 3081
rect 3311 3060 3315 3091
rect 3409 3067 3566 3071
rect 3409 3060 3413 3067
rect 3311 3056 3413 3060
rect 3562 3050 3566 3067
rect 3597 3064 3601 3173
rect 3622 3085 3626 3151
rect 3246 2507 3250 2784
rect 3622 2607 3626 3074
rect 3643 3050 3647 3051
rect 3622 2500 3626 2573
rect 3248 2341 3252 2496
rect 3241 1936 3309 1940
rect 3241 1915 3245 1936
rect 3248 1763 3252 1925
rect 3305 1904 3309 1936
rect 3409 1911 3565 1915
rect 3409 1904 3413 1911
rect 3305 1900 3413 1904
rect 3561 1894 3565 1911
rect 3597 1908 3601 2017
rect 3622 1929 3626 1995
rect 3246 1351 3250 1628
rect 3622 1451 3626 1918
rect 3622 1344 3626 1417
rect 3650 1405 3658 3508
rect 3661 3057 3665 3631
rect 3661 2479 3665 3053
rect 3661 1901 3665 2475
rect 3668 2927 3672 3501
rect 3668 2349 3672 2923
rect 3668 1771 3672 2345
rect 3402 1272 3406 1340
rect 3499 1272 3503 1340
rect 3650 1040 3658 1398
rect 2642 1000 2654 1028
rect 2708 1027 2716 1028
rect 3179 1027 3187 1028
rect 2602 996 2698 1000
rect 2620 994 2634 996
use DMUX  DMUX_0
timestamp 1414996929
transform 1 0 1254 0 1 3642
box -19 3 78 111
use MUX2X1  MUX2X1_5
timestamp 1414990262
transform 1 0 1816 0 1 3648
box -5 -3 53 105
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 1858 0 1 3648
box -9 -3 26 105
use OR2X1  OR2X1_0
timestamp 1053022145
transform 1 0 2243 0 1 3648
box -8 -3 40 105
use DMUX  DMUX_2
timestamp 1414996929
transform 1 0 2667 0 1 3642
box -19 3 78 111
use MUX2X1  MUX2X1_6
timestamp 1414990262
transform 1 0 2758 0 1 3648
box -5 -3 53 105
use INVX1  INVX1_1
timestamp 1053022145
transform 1 0 2800 0 1 3648
box -9 -3 26 105
use DMUX  DMUX_4
timestamp 1414996929
transform 1 0 3138 0 1 3642
box -19 3 78 111
use DMUX  DMUX_1
timestamp 1414996929
transform 1 0 1255 0 1 3526
box -19 3 78 111
use MUX2X1  MUX2X1_4
timestamp 1414990262
transform 1 0 1228 0 1 2659
box -5 -3 53 105
use DMUX  DMUX_3
timestamp 1414996929
transform 1 0 1238 0 1 1995
box -19 3 78 111
use MUX2X1  MUX2X1_0
timestamp 1414990262
transform 1 0 1238 0 1 1459
box -5 -3 53 105
use MUX2X1  MUX2X1_7
timestamp 1414990262
transform 1 0 3702 0 1 3272
box -5 -3 53 105
use DMUX  DMUX_5
timestamp 1414996929
transform 1 0 3708 0 1 2624
box -19 3 78 111
use MUX2X1  MUX2X1_8
timestamp 1414990262
transform 1 0 3700 0 1 2110
box -5 -3 53 105
use DMUX  DMUX_6
timestamp 1414996929
transform 1 0 3694 0 1 1435
box -19 3 78 111
use PLU  PLU_0
array 0 4 471 0 3 578
timestamp 1414992301
transform 1 0 1326 0 1 1377
box -9 -40 462 538
use MUX2X1  MUX2X1_1
timestamp 1414990262
transform 1 0 1363 0 1 1240
box -5 -3 53 105
use DMUX  DMUX_7
timestamp 1414996929
transform 1 0 2028 0 1 1211
box -19 3 78 111
use MUX2X1  MUX2X1_2
timestamp 1414990262
transform 1 0 2335 0 1 1227
box -5 -3 53 105
use DMUX  DMUX_8
timestamp 1414996929
transform 1 0 2982 0 1 1214
box -19 3 78 111
use MUX2X1  MUX2X1_3
timestamp 1414990262
transform 1 0 3286 0 1 1228
box -5 -3 53 105
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1415033039
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
