* SPICE 3f5 Level 8, Star-HSPICE Level 49, UTMOST Level 8

* DATE: Aug 13/03
* LOT: T36S                  WAF: 1101
* Temperature_parameters=Default
.MODEL nfet NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6461285
+K1      = 0.9152455      K2      = -0.105898      K3      = 26.1007653
+K3B     = -8.3258109     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 3.7861788      DVT1    = 0.3717718      DVT2    = -0.0830195
+U0      = 442.2002499    UA      = 1E-13          UB      = 1.185519E-18
+UC      = 6.470959E-12   VSAT    = 1.727533E5     A0      = 0.6072333
+AGS     = 0.1377586      B0      = 2.667083E-6    B1      = 5E-6
+KETA    = -2.897119E-3   A1      = 3.028408E-4    A2      = 0.345619
+RDSW    = 1.077249E3     PRWG    = 0.1399237      PRWB    = 0.0595509
+WR      = 1              WINT    = 2.208544E-7    LINT    = 4.960111E-8
+XL      = 1E-7           XW      = 0              DWG     = -1.893724E-9
+DWB     = 5.47692E-8     VOFF    = 0              NFACTOR = 0.472999
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 2.181479E-3    ETAB    = -6.299339E-4
+DSUB    = 0.0689754      PCLM    = 2.4881989      PDIBLC1 = 0.9941032
+PDIBLC2 = 2.298113E-3    PDIBLCB = -0.0180618     DROUT   = 0.8838803
+PSCBE1  = 6.445443E8     PSCBE2  = 2.598335E-4    PVAG    = 0
+DELTA   = 0.01           RSH     = 81.8           MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.01E-10       CGSO    = 2.01E-10       CGBO    = 1E-9
+CJ      = 4.227962E-4    PB      = 0.9113851      MJ      = 0.4296861
+CJSW    = 2.925306E-10   PBSW    = 0.8            MJSW    = 0.170165
+CJSWG   = 1.64E-10       PBSWG   = 0.8            MJSWG   = 0.170165
+CF      = 0              PVTH0   = 0.1375778      PRDSW   = -174.8924404
+PK2     = -0.0194887     WKETA   = -0.0237035     LKETA   = 0.0205439       )
*
.MODEL pfet PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9213369
+K1      = 0.5309886      K2      = 0.0157077      K3      = 3.9841467
+K3B     = -0.8977975     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.8313335      DVT1    = 0.4250351      DVT2    = -0.055987
+U0      = 209.2163727    UA      = 2.878347E-9    UB      = 1.397451E-21
+UC      = -6.27575E-11   VSAT    = 2E5            A0      = 0.9102666
+AGS     = 0.1449591      B0      = 1.211218E-6    B1      = 5E-6
+KETA    = -1.616658E-3   A1      = 0              A2      = 0.3
+RDSW    = 2.088968E3     PRWG    = 2.930817E-4    PRWB    = -0.0963307
+WR      = 1              WINT    = 3.279186E-7    LINT    = 6.251424E-8
+XL      = 1E-7           XW      = 0              DWG     = -2.846864E-8
+DWB     = 1.437983E-8    VOFF    = -0.0130604     NFACTOR = 1.0218439
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.1086822      ETAB    = -0.0677706
+DSUB    = 0.8682467      PCLM    = 2.168708       PDIBLC1 = 0.112826
+PDIBLC2 = 3.525757E-3    PDIBLCB = -0.059791      DROUT   = 0.3016682
+PSCBE1  = 5.091678E9     PSCBE2  = 5E-10          PVAG    = 0.0256592
+DELTA   = 0.01           RSH     = 102            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.62E-10       CGSO    = 2.62E-10       CGBO    = 1E-9
+CJ      = 7.247826E-4    PB      = 0.9541788      MJ      = 0.4958349
+CJSW    = 2.613323E-10   PBSW    = 0.99           MJSW    = 0.2516611
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.2516611
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 3.391823E-3    LKETA   = -8.97011E-3     )
*
